module Instr_Mem #(parameter PROG_CTR_WID = 10) (
	input clk,	input [PROG_CTR_WID-1:0] prog_ctr,
	output reg [15:0] instr_mem_out
);
always @(posedge clk) begin
	case (prog_ctr)
		10'h000: instr_mem_out <= 16'h963F;
		10'h001: instr_mem_out <= 16'h970D;
		10'h002: instr_mem_out <= 16'h0000;
		10'h003: instr_mem_out <= 16'h0000;
		10'h004: instr_mem_out <= 16'hD601;
		10'h005: instr_mem_out <= 16'hD701;
		10'h006: instr_mem_out <= 16'h0000;
		10'h007: instr_mem_out <= 16'h0000;
		10'h008: instr_mem_out <= 16'h0000;
		10'h009: instr_mem_out <= 16'hD601;
		10'h00A: instr_mem_out <= 16'hD701;
		10'h00B: instr_mem_out <= 16'h0000;
		10'h00C: instr_mem_out <= 16'h0000;
		10'h00D: instr_mem_out <= 16'h0000;
		10'h00E: instr_mem_out <= 16'hD601;
		10'h00F: instr_mem_out <= 16'hD701;
		10'h010: instr_mem_out <= 16'h0000;
		10'h011: instr_mem_out <= 16'h0000;
		10'h012: instr_mem_out <= 16'h0000;
		10'h013: instr_mem_out <= 16'hD601;
		10'h014: instr_mem_out <= 16'hD701;
		10'h015: instr_mem_out <= 16'h0000;
		10'h016: instr_mem_out <= 16'h0000;
		10'h017: instr_mem_out <= 16'h0000;
		10'h018: instr_mem_out <= 16'hD601;
		10'h019: instr_mem_out <= 16'hD701;
		10'h01A: instr_mem_out <= 16'h0000;
		10'h01B: instr_mem_out <= 16'h0000;
		10'h01C: instr_mem_out <= 16'h0000;
		10'h01D: instr_mem_out <= 16'hD601;
		10'h01E: instr_mem_out <= 16'hD701;
		10'h01F: instr_mem_out <= 16'h0000;
		10'h020: instr_mem_out <= 16'h0000;
		10'h021: instr_mem_out <= 16'h0000;
		10'h022: instr_mem_out <= 16'hD601;
		10'h023: instr_mem_out <= 16'hD701;
		10'h024: instr_mem_out <= 16'h0000;
		10'h025: instr_mem_out <= 16'h0000;
		10'h026: instr_mem_out <= 16'h0000;
		10'h027: instr_mem_out <= 16'hD601;
		10'h028: instr_mem_out <= 16'hD701;
		10'h029: instr_mem_out <= 16'h0000;
		10'h02A: instr_mem_out <= 16'h0000;
		10'h02B: instr_mem_out <= 16'h0000;
		10'h02C: instr_mem_out <= 16'hD601;
		10'h02D: instr_mem_out <= 16'hD701;
		10'h02E: instr_mem_out <= 16'h0000;
		10'h02F: instr_mem_out <= 16'h0000;
		10'h030: instr_mem_out <= 16'h0000;
		10'h031: instr_mem_out <= 16'hD601;
		10'h032: instr_mem_out <= 16'hD701;
		10'h033: instr_mem_out <= 16'h0000;
		10'h034: instr_mem_out <= 16'h0000;
		10'h035: instr_mem_out <= 16'h0000;
		10'h036: instr_mem_out <= 16'hD601;
		10'h037: instr_mem_out <= 16'hD701;
		10'h038: instr_mem_out <= 16'h0000;
		10'h039: instr_mem_out <= 16'h0000;
		10'h03A: instr_mem_out <= 16'h0000;
		10'h03B: instr_mem_out <= 16'hD601;
		10'h03C: instr_mem_out <= 16'hD701;
		10'h03D: instr_mem_out <= 16'h0000;
		10'h03E: instr_mem_out <= 16'h0000;
		10'h03F: instr_mem_out <= 16'h0000;
		10'h040: instr_mem_out <= 16'hD601;
		10'h041: instr_mem_out <= 16'hD701;
		10'h042: instr_mem_out <= 16'h0000;
		10'h043: instr_mem_out <= 16'h0000;
		10'h044: instr_mem_out <= 16'h0000;
		10'h045: instr_mem_out <= 16'h9011;
		10'h046: instr_mem_out <= 16'h9122;
		10'h047: instr_mem_out <= 16'h9810;
		10'h048: instr_mem_out <= 16'hA101;
		10'h049: instr_mem_out <= 16'hAA11;
		10'h04A: instr_mem_out <= 16'hBA08;
		10'h04B: instr_mem_out <= 16'hD201;
		10'h04C: instr_mem_out <= 16'hC208;
		10'h04D: instr_mem_out <= 16'hD201;
		10'h04E: instr_mem_out <= 16'hBA09;
		10'h04F: instr_mem_out <= 16'hD201;
		10'h050: instr_mem_out <= 16'hC209;
		10'h051: instr_mem_out <= 16'hD201;
		10'h052: instr_mem_out <= 16'hBA0A;
		10'h053: instr_mem_out <= 16'hD201;
		10'h054: instr_mem_out <= 16'hC20A;
		10'h055: instr_mem_out <= 16'hD201;
		10'h056: instr_mem_out <= 16'h9001;
		10'h057: instr_mem_out <= 16'h9101;
		10'h058: instr_mem_out <= 16'h9281;
		10'h059: instr_mem_out <= 16'h96FF;
		10'h05A: instr_mem_out <= 16'hD601;
		10'h05B: instr_mem_out <= 16'hD601;
		10'h05C: instr_mem_out <= 16'hD601;
		10'h05D: instr_mem_out <= 16'hD601;
		10'h05E: instr_mem_out <= 16'hD601;
		10'h05F: instr_mem_out <= 16'hD601;
		10'h060: instr_mem_out <= 16'hD601;
		10'h061: instr_mem_out <= 16'hD601;
		10'h062: instr_mem_out <= 16'hD601;
		10'h063: instr_mem_out <= 16'hD601;
		10'h064: instr_mem_out <= 16'hD601;
		10'h065: instr_mem_out <= 16'hA800;
		10'h066: instr_mem_out <= 16'hBB08;
		10'h067: instr_mem_out <= 16'hC408;
		10'h068: instr_mem_out <= 16'hD301;
		10'h069: instr_mem_out <= 16'hD401;
		10'h06A: instr_mem_out <= 16'h0810;
		10'h06B: instr_mem_out <= 16'h6820;
		10'h06C: instr_mem_out <= 16'h8073;
		10'h06D: instr_mem_out <= 16'hDD03;
		10'h06E: instr_mem_out <= 16'h0000;
		10'h06F: instr_mem_out <= 16'h6865;
		10'h070: instr_mem_out <= 16'h806D;
		10'h071: instr_mem_out <= 16'h3865;
		10'h072: instr_mem_out <= 16'h0000;
		10'h073: instr_mem_out <= 16'hDD02;
		10'h074: instr_mem_out <= 16'h0000;
		10'h075: instr_mem_out <= 16'h6865;
		10'h076: instr_mem_out <= 16'h7872;
		10'h077: instr_mem_out <= 16'hDD03;
		10'h078: instr_mem_out <= 16'h0000;
		10'h079: instr_mem_out <= 16'h6865;
		10'h07A: instr_mem_out <= 16'h8077;
		10'h07B: instr_mem_out <= 16'hDD01;
		10'h07C: instr_mem_out <= 16'h0000;
		10'h07D: instr_mem_out <= 16'hD501;
		10'h07E: instr_mem_out <= 16'h3873;
		10'h07F: instr_mem_out <= 16'h0000;
		10'h080: instr_mem_out <= 16'h0000;
		10'h081: instr_mem_out <= 16'h0000;
		10'h082: instr_mem_out <= 16'h0000;
		10'h083: instr_mem_out <= 16'h0000;
		10'h084: instr_mem_out <= 16'h0000;
		10'h085: instr_mem_out <= 16'h0000;
		10'h086: instr_mem_out <= 16'h0000;
		10'h087: instr_mem_out <= 16'h0000;
		10'h088: instr_mem_out <= 16'h0000;
		10'h089: instr_mem_out <= 16'h0000;
		10'h08A: instr_mem_out <= 16'h0000;
		10'h08B: instr_mem_out <= 16'h0000;
		10'h08C: instr_mem_out <= 16'h0000;
		10'h08D: instr_mem_out <= 16'h0000;
		10'h08E: instr_mem_out <= 16'h0000;
		10'h08F: instr_mem_out <= 16'h0000;
		10'h090: instr_mem_out <= 16'h0000;
		10'h091: instr_mem_out <= 16'h0000;
		10'h092: instr_mem_out <= 16'h0000;
		10'h093: instr_mem_out <= 16'h0000;
		10'h094: instr_mem_out <= 16'h0000;
		10'h095: instr_mem_out <= 16'h0000;
		10'h096: instr_mem_out <= 16'h0000;
		10'h097: instr_mem_out <= 16'h0000;
		10'h098: instr_mem_out <= 16'h0000;
		10'h099: instr_mem_out <= 16'h0000;
		10'h09A: instr_mem_out <= 16'h0000;
		10'h09B: instr_mem_out <= 16'h0000;
		10'h09C: instr_mem_out <= 16'h0000;
		10'h09D: instr_mem_out <= 16'h0000;
		10'h09E: instr_mem_out <= 16'h0000;
		10'h09F: instr_mem_out <= 16'h0000;
		10'h0A0: instr_mem_out <= 16'h0000;
		10'h0A1: instr_mem_out <= 16'h0000;
		10'h0A2: instr_mem_out <= 16'h0000;
		10'h0A3: instr_mem_out <= 16'h0000;
		10'h0A4: instr_mem_out <= 16'h0000;
		10'h0A5: instr_mem_out <= 16'h0000;
		10'h0A6: instr_mem_out <= 16'h0000;
		10'h0A7: instr_mem_out <= 16'h0000;
		10'h0A8: instr_mem_out <= 16'h0000;
		10'h0A9: instr_mem_out <= 16'h0000;
		10'h0AA: instr_mem_out <= 16'h0000;
		10'h0AB: instr_mem_out <= 16'h0000;
		10'h0AC: instr_mem_out <= 16'h0000;
		10'h0AD: instr_mem_out <= 16'h0000;
		10'h0AE: instr_mem_out <= 16'h0000;
		10'h0AF: instr_mem_out <= 16'h0000;
		10'h0B0: instr_mem_out <= 16'h0000;
		10'h0B1: instr_mem_out <= 16'h0000;
		10'h0B2: instr_mem_out <= 16'h0000;
		10'h0B3: instr_mem_out <= 16'h0000;
		10'h0B4: instr_mem_out <= 16'h0000;
		10'h0B5: instr_mem_out <= 16'h0000;
		10'h0B6: instr_mem_out <= 16'h0000;
		10'h0B7: instr_mem_out <= 16'h0000;
		10'h0B8: instr_mem_out <= 16'h0000;
		10'h0B9: instr_mem_out <= 16'h0000;
		10'h0BA: instr_mem_out <= 16'h0000;
		10'h0BB: instr_mem_out <= 16'h0000;
		10'h0BC: instr_mem_out <= 16'h0000;
		10'h0BD: instr_mem_out <= 16'h0000;
		10'h0BE: instr_mem_out <= 16'h0000;
		10'h0BF: instr_mem_out <= 16'h0000;
		10'h0C0: instr_mem_out <= 16'h0000;
		10'h0C1: instr_mem_out <= 16'h0000;
		10'h0C2: instr_mem_out <= 16'h0000;
		10'h0C3: instr_mem_out <= 16'h0000;
		10'h0C4: instr_mem_out <= 16'h0000;
		10'h0C5: instr_mem_out <= 16'h0000;
		10'h0C6: instr_mem_out <= 16'h0000;
		10'h0C7: instr_mem_out <= 16'h0000;
		10'h0C8: instr_mem_out <= 16'h0000;
		10'h0C9: instr_mem_out <= 16'h0000;
		10'h0CA: instr_mem_out <= 16'h0000;
		10'h0CB: instr_mem_out <= 16'h0000;
		10'h0CC: instr_mem_out <= 16'h0000;
		10'h0CD: instr_mem_out <= 16'h0000;
		10'h0CE: instr_mem_out <= 16'h0000;
		10'h0CF: instr_mem_out <= 16'h0000;
		10'h0D0: instr_mem_out <= 16'h0000;
		10'h0D1: instr_mem_out <= 16'h0000;
		10'h0D2: instr_mem_out <= 16'h0000;
		10'h0D3: instr_mem_out <= 16'h0000;
		10'h0D4: instr_mem_out <= 16'h0000;
		10'h0D5: instr_mem_out <= 16'h0000;
		10'h0D6: instr_mem_out <= 16'h0000;
		10'h0D7: instr_mem_out <= 16'h0000;
		10'h0D8: instr_mem_out <= 16'h0000;
		10'h0D9: instr_mem_out <= 16'h0000;
		10'h0DA: instr_mem_out <= 16'h0000;
		10'h0DB: instr_mem_out <= 16'h0000;
		10'h0DC: instr_mem_out <= 16'h0000;
		10'h0DD: instr_mem_out <= 16'h0000;
		10'h0DE: instr_mem_out <= 16'h0000;
		10'h0DF: instr_mem_out <= 16'h0000;
		10'h0E0: instr_mem_out <= 16'h0000;
		10'h0E1: instr_mem_out <= 16'h0000;
		10'h0E2: instr_mem_out <= 16'h0000;
		10'h0E3: instr_mem_out <= 16'h0000;
		10'h0E4: instr_mem_out <= 16'h0000;
		10'h0E5: instr_mem_out <= 16'h0000;
		10'h0E6: instr_mem_out <= 16'h0000;
		10'h0E7: instr_mem_out <= 16'h0000;
		10'h0E8: instr_mem_out <= 16'h0000;
		10'h0E9: instr_mem_out <= 16'h0000;
		10'h0EA: instr_mem_out <= 16'h0000;
		10'h0EB: instr_mem_out <= 16'h0000;
		10'h0EC: instr_mem_out <= 16'h0000;
		10'h0ED: instr_mem_out <= 16'h0000;
		10'h0EE: instr_mem_out <= 16'h0000;
		10'h0EF: instr_mem_out <= 16'h0000;
		10'h0F0: instr_mem_out <= 16'h0000;
		10'h0F1: instr_mem_out <= 16'h0000;
		10'h0F2: instr_mem_out <= 16'h0000;
		10'h0F3: instr_mem_out <= 16'h0000;
		10'h0F4: instr_mem_out <= 16'h0000;
		10'h0F5: instr_mem_out <= 16'h0000;
		10'h0F6: instr_mem_out <= 16'h0000;
		10'h0F7: instr_mem_out <= 16'h0000;
		10'h0F8: instr_mem_out <= 16'h0000;
		10'h0F9: instr_mem_out <= 16'h0000;
		10'h0FA: instr_mem_out <= 16'h0000;
		10'h0FB: instr_mem_out <= 16'h0000;
		10'h0FC: instr_mem_out <= 16'h0000;
		10'h0FD: instr_mem_out <= 16'h0000;
		10'h0FE: instr_mem_out <= 16'h0000;
		10'h0FF: instr_mem_out <= 16'h0000;
		10'h100: instr_mem_out <= 16'h0000;
		10'h101: instr_mem_out <= 16'h0000;
		10'h102: instr_mem_out <= 16'h0000;
		10'h103: instr_mem_out <= 16'h0000;
		10'h104: instr_mem_out <= 16'h0000;
		10'h105: instr_mem_out <= 16'h0000;
		10'h106: instr_mem_out <= 16'h0000;
		10'h107: instr_mem_out <= 16'h0000;
		10'h108: instr_mem_out <= 16'h0000;
		10'h109: instr_mem_out <= 16'h0000;
		10'h10A: instr_mem_out <= 16'h0000;
		10'h10B: instr_mem_out <= 16'h0000;
		10'h10C: instr_mem_out <= 16'h0000;
		10'h10D: instr_mem_out <= 16'h0000;
		10'h10E: instr_mem_out <= 16'h0000;
		10'h10F: instr_mem_out <= 16'h0000;
		10'h110: instr_mem_out <= 16'h0000;
		10'h111: instr_mem_out <= 16'h0000;
		10'h112: instr_mem_out <= 16'h0000;
		10'h113: instr_mem_out <= 16'h0000;
		10'h114: instr_mem_out <= 16'h0000;
		10'h115: instr_mem_out <= 16'h0000;
		10'h116: instr_mem_out <= 16'h0000;
		10'h117: instr_mem_out <= 16'h0000;
		10'h118: instr_mem_out <= 16'h0000;
		10'h119: instr_mem_out <= 16'h0000;
		10'h11A: instr_mem_out <= 16'h0000;
		10'h11B: instr_mem_out <= 16'h0000;
		10'h11C: instr_mem_out <= 16'h0000;
		10'h11D: instr_mem_out <= 16'h0000;
		10'h11E: instr_mem_out <= 16'h0000;
		10'h11F: instr_mem_out <= 16'h0000;
		10'h120: instr_mem_out <= 16'h0000;
		10'h121: instr_mem_out <= 16'h0000;
		10'h122: instr_mem_out <= 16'h0000;
		10'h123: instr_mem_out <= 16'h0000;
		10'h124: instr_mem_out <= 16'h0000;
		10'h125: instr_mem_out <= 16'h0000;
		10'h126: instr_mem_out <= 16'h0000;
		10'h127: instr_mem_out <= 16'h0000;
		10'h128: instr_mem_out <= 16'h0000;
		10'h129: instr_mem_out <= 16'h0000;
		10'h12A: instr_mem_out <= 16'h0000;
		10'h12B: instr_mem_out <= 16'h0000;
		10'h12C: instr_mem_out <= 16'h0000;
		10'h12D: instr_mem_out <= 16'h0000;
		10'h12E: instr_mem_out <= 16'h0000;
		10'h12F: instr_mem_out <= 16'h0000;
		10'h130: instr_mem_out <= 16'h0000;
		10'h131: instr_mem_out <= 16'h0000;
		10'h132: instr_mem_out <= 16'h0000;
		10'h133: instr_mem_out <= 16'h0000;
		10'h134: instr_mem_out <= 16'h0000;
		10'h135: instr_mem_out <= 16'h0000;
		10'h136: instr_mem_out <= 16'h0000;
		10'h137: instr_mem_out <= 16'h0000;
		10'h138: instr_mem_out <= 16'h0000;
		10'h139: instr_mem_out <= 16'h0000;
		10'h13A: instr_mem_out <= 16'h0000;
		10'h13B: instr_mem_out <= 16'h0000;
		10'h13C: instr_mem_out <= 16'h0000;
		10'h13D: instr_mem_out <= 16'h0000;
		10'h13E: instr_mem_out <= 16'h0000;
		10'h13F: instr_mem_out <= 16'h0000;
		10'h140: instr_mem_out <= 16'h0000;
		10'h141: instr_mem_out <= 16'h0000;
		10'h142: instr_mem_out <= 16'h0000;
		10'h143: instr_mem_out <= 16'h0000;
		10'h144: instr_mem_out <= 16'h0000;
		10'h145: instr_mem_out <= 16'h0000;
		10'h146: instr_mem_out <= 16'h0000;
		10'h147: instr_mem_out <= 16'h0000;
		10'h148: instr_mem_out <= 16'h0000;
		10'h149: instr_mem_out <= 16'h0000;
		10'h14A: instr_mem_out <= 16'h0000;
		10'h14B: instr_mem_out <= 16'h0000;
		10'h14C: instr_mem_out <= 16'h0000;
		10'h14D: instr_mem_out <= 16'h0000;
		10'h14E: instr_mem_out <= 16'h0000;
		10'h14F: instr_mem_out <= 16'h0000;
		10'h150: instr_mem_out <= 16'h0000;
		10'h151: instr_mem_out <= 16'h0000;
		10'h152: instr_mem_out <= 16'h0000;
		10'h153: instr_mem_out <= 16'h0000;
		10'h154: instr_mem_out <= 16'h0000;
		10'h155: instr_mem_out <= 16'h0000;
		10'h156: instr_mem_out <= 16'h0000;
		10'h157: instr_mem_out <= 16'h0000;
		10'h158: instr_mem_out <= 16'h0000;
		10'h159: instr_mem_out <= 16'h0000;
		10'h15A: instr_mem_out <= 16'h0000;
		10'h15B: instr_mem_out <= 16'h0000;
		10'h15C: instr_mem_out <= 16'h0000;
		10'h15D: instr_mem_out <= 16'h0000;
		10'h15E: instr_mem_out <= 16'h0000;
		10'h15F: instr_mem_out <= 16'h0000;
		10'h160: instr_mem_out <= 16'h0000;
		10'h161: instr_mem_out <= 16'h0000;
		10'h162: instr_mem_out <= 16'h0000;
		10'h163: instr_mem_out <= 16'h0000;
		10'h164: instr_mem_out <= 16'h0000;
		10'h165: instr_mem_out <= 16'h0000;
		10'h166: instr_mem_out <= 16'h0000;
		10'h167: instr_mem_out <= 16'h0000;
		10'h168: instr_mem_out <= 16'h0000;
		10'h169: instr_mem_out <= 16'h0000;
		10'h16A: instr_mem_out <= 16'h0000;
		10'h16B: instr_mem_out <= 16'h0000;
		10'h16C: instr_mem_out <= 16'h0000;
		10'h16D: instr_mem_out <= 16'h0000;
		10'h16E: instr_mem_out <= 16'h0000;
		10'h16F: instr_mem_out <= 16'h0000;
		10'h170: instr_mem_out <= 16'h0000;
		10'h171: instr_mem_out <= 16'h0000;
		10'h172: instr_mem_out <= 16'h0000;
		10'h173: instr_mem_out <= 16'h0000;
		10'h174: instr_mem_out <= 16'h0000;
		10'h175: instr_mem_out <= 16'h0000;
		10'h176: instr_mem_out <= 16'h0000;
		10'h177: instr_mem_out <= 16'h0000;
		10'h178: instr_mem_out <= 16'h0000;
		10'h179: instr_mem_out <= 16'h0000;
		10'h17A: instr_mem_out <= 16'h0000;
		10'h17B: instr_mem_out <= 16'h0000;
		10'h17C: instr_mem_out <= 16'h0000;
		10'h17D: instr_mem_out <= 16'h0000;
		10'h17E: instr_mem_out <= 16'h0000;
		10'h17F: instr_mem_out <= 16'h0000;
		10'h180: instr_mem_out <= 16'h0000;
		10'h181: instr_mem_out <= 16'h0000;
		10'h182: instr_mem_out <= 16'h0000;
		10'h183: instr_mem_out <= 16'h0000;
		10'h184: instr_mem_out <= 16'h0000;
		10'h185: instr_mem_out <= 16'h0000;
		10'h186: instr_mem_out <= 16'h0000;
		10'h187: instr_mem_out <= 16'h0000;
		10'h188: instr_mem_out <= 16'h0000;
		10'h189: instr_mem_out <= 16'h0000;
		10'h18A: instr_mem_out <= 16'h0000;
		10'h18B: instr_mem_out <= 16'h0000;
		10'h18C: instr_mem_out <= 16'h0000;
		10'h18D: instr_mem_out <= 16'h0000;
		10'h18E: instr_mem_out <= 16'h0000;
		10'h18F: instr_mem_out <= 16'h0000;
		10'h190: instr_mem_out <= 16'h0000;
		10'h191: instr_mem_out <= 16'h0000;
		10'h192: instr_mem_out <= 16'h0000;
		10'h193: instr_mem_out <= 16'h0000;
		10'h194: instr_mem_out <= 16'h0000;
		10'h195: instr_mem_out <= 16'h0000;
		10'h196: instr_mem_out <= 16'h0000;
		10'h197: instr_mem_out <= 16'h0000;
		10'h198: instr_mem_out <= 16'h0000;
		10'h199: instr_mem_out <= 16'h0000;
		10'h19A: instr_mem_out <= 16'h0000;
		10'h19B: instr_mem_out <= 16'h0000;
		10'h19C: instr_mem_out <= 16'h0000;
		10'h19D: instr_mem_out <= 16'h0000;
		10'h19E: instr_mem_out <= 16'h0000;
		10'h19F: instr_mem_out <= 16'h0000;
		10'h1A0: instr_mem_out <= 16'h0000;
		10'h1A1: instr_mem_out <= 16'h0000;
		10'h1A2: instr_mem_out <= 16'h0000;
		10'h1A3: instr_mem_out <= 16'h0000;
		10'h1A4: instr_mem_out <= 16'h0000;
		10'h1A5: instr_mem_out <= 16'h0000;
		10'h1A6: instr_mem_out <= 16'h0000;
		10'h1A7: instr_mem_out <= 16'h0000;
		10'h1A8: instr_mem_out <= 16'h0000;
		10'h1A9: instr_mem_out <= 16'h0000;
		10'h1AA: instr_mem_out <= 16'h0000;
		10'h1AB: instr_mem_out <= 16'h0000;
		10'h1AC: instr_mem_out <= 16'h0000;
		10'h1AD: instr_mem_out <= 16'h0000;
		10'h1AE: instr_mem_out <= 16'h0000;
		10'h1AF: instr_mem_out <= 16'h0000;
		10'h1B0: instr_mem_out <= 16'h0000;
		10'h1B1: instr_mem_out <= 16'h0000;
		10'h1B2: instr_mem_out <= 16'h0000;
		10'h1B3: instr_mem_out <= 16'h0000;
		10'h1B4: instr_mem_out <= 16'h0000;
		10'h1B5: instr_mem_out <= 16'h0000;
		10'h1B6: instr_mem_out <= 16'h0000;
		10'h1B7: instr_mem_out <= 16'h0000;
		10'h1B8: instr_mem_out <= 16'h0000;
		10'h1B9: instr_mem_out <= 16'h0000;
		10'h1BA: instr_mem_out <= 16'h0000;
		10'h1BB: instr_mem_out <= 16'h0000;
		10'h1BC: instr_mem_out <= 16'h0000;
		10'h1BD: instr_mem_out <= 16'h0000;
		10'h1BE: instr_mem_out <= 16'h0000;
		10'h1BF: instr_mem_out <= 16'h0000;
		10'h1C0: instr_mem_out <= 16'h0000;
		10'h1C1: instr_mem_out <= 16'h0000;
		10'h1C2: instr_mem_out <= 16'h0000;
		10'h1C3: instr_mem_out <= 16'h0000;
		10'h1C4: instr_mem_out <= 16'h0000;
		10'h1C5: instr_mem_out <= 16'h0000;
		10'h1C6: instr_mem_out <= 16'h0000;
		10'h1C7: instr_mem_out <= 16'h0000;
		10'h1C8: instr_mem_out <= 16'h0000;
		10'h1C9: instr_mem_out <= 16'h0000;
		10'h1CA: instr_mem_out <= 16'h0000;
		10'h1CB: instr_mem_out <= 16'h0000;
		10'h1CC: instr_mem_out <= 16'h0000;
		10'h1CD: instr_mem_out <= 16'h0000;
		10'h1CE: instr_mem_out <= 16'h0000;
		10'h1CF: instr_mem_out <= 16'h0000;
		10'h1D0: instr_mem_out <= 16'h0000;
		10'h1D1: instr_mem_out <= 16'h0000;
		10'h1D2: instr_mem_out <= 16'h0000;
		10'h1D3: instr_mem_out <= 16'h0000;
		10'h1D4: instr_mem_out <= 16'h0000;
		10'h1D5: instr_mem_out <= 16'h0000;
		10'h1D6: instr_mem_out <= 16'h0000;
		10'h1D7: instr_mem_out <= 16'h0000;
		10'h1D8: instr_mem_out <= 16'h0000;
		10'h1D9: instr_mem_out <= 16'h0000;
		10'h1DA: instr_mem_out <= 16'h0000;
		10'h1DB: instr_mem_out <= 16'h0000;
		10'h1DC: instr_mem_out <= 16'h0000;
		10'h1DD: instr_mem_out <= 16'h0000;
		10'h1DE: instr_mem_out <= 16'h0000;
		10'h1DF: instr_mem_out <= 16'h0000;
		10'h1E0: instr_mem_out <= 16'h0000;
		10'h1E1: instr_mem_out <= 16'h0000;
		10'h1E2: instr_mem_out <= 16'h0000;
		10'h1E3: instr_mem_out <= 16'h0000;
		10'h1E4: instr_mem_out <= 16'h0000;
		10'h1E5: instr_mem_out <= 16'h0000;
		10'h1E6: instr_mem_out <= 16'h0000;
		10'h1E7: instr_mem_out <= 16'h0000;
		10'h1E8: instr_mem_out <= 16'h0000;
		10'h1E9: instr_mem_out <= 16'h0000;
		10'h1EA: instr_mem_out <= 16'h0000;
		10'h1EB: instr_mem_out <= 16'h0000;
		10'h1EC: instr_mem_out <= 16'h0000;
		10'h1ED: instr_mem_out <= 16'h0000;
		10'h1EE: instr_mem_out <= 16'h0000;
		10'h1EF: instr_mem_out <= 16'h0000;
		10'h1F0: instr_mem_out <= 16'h0000;
		10'h1F1: instr_mem_out <= 16'h0000;
		10'h1F2: instr_mem_out <= 16'h0000;
		10'h1F3: instr_mem_out <= 16'h0000;
		10'h1F4: instr_mem_out <= 16'h0000;
		10'h1F5: instr_mem_out <= 16'h0000;
		10'h1F6: instr_mem_out <= 16'h0000;
		10'h1F7: instr_mem_out <= 16'h0000;
		10'h1F8: instr_mem_out <= 16'h0000;
		10'h1F9: instr_mem_out <= 16'h0000;
		10'h1FA: instr_mem_out <= 16'h0000;
		10'h1FB: instr_mem_out <= 16'h0000;
		10'h1FC: instr_mem_out <= 16'h0000;
		10'h1FD: instr_mem_out <= 16'h0000;
		10'h1FE: instr_mem_out <= 16'h0000;
		10'h1FF: instr_mem_out <= 16'h0000;
		10'h200: instr_mem_out <= 16'h0000;
		10'h201: instr_mem_out <= 16'h0000;
		10'h202: instr_mem_out <= 16'h0000;
		10'h203: instr_mem_out <= 16'h0000;
		10'h204: instr_mem_out <= 16'h0000;
		10'h205: instr_mem_out <= 16'h0000;
		10'h206: instr_mem_out <= 16'h0000;
		10'h207: instr_mem_out <= 16'h0000;
		10'h208: instr_mem_out <= 16'h0000;
		10'h209: instr_mem_out <= 16'h0000;
		10'h20A: instr_mem_out <= 16'h0000;
		10'h20B: instr_mem_out <= 16'h0000;
		10'h20C: instr_mem_out <= 16'h0000;
		10'h20D: instr_mem_out <= 16'h0000;
		10'h20E: instr_mem_out <= 16'h0000;
		10'h20F: instr_mem_out <= 16'h0000;
		10'h210: instr_mem_out <= 16'h0000;
		10'h211: instr_mem_out <= 16'h0000;
		10'h212: instr_mem_out <= 16'h0000;
		10'h213: instr_mem_out <= 16'h0000;
		10'h214: instr_mem_out <= 16'h0000;
		10'h215: instr_mem_out <= 16'h0000;
		10'h216: instr_mem_out <= 16'h0000;
		10'h217: instr_mem_out <= 16'h0000;
		10'h218: instr_mem_out <= 16'h0000;
		10'h219: instr_mem_out <= 16'h0000;
		10'h21A: instr_mem_out <= 16'h0000;
		10'h21B: instr_mem_out <= 16'h0000;
		10'h21C: instr_mem_out <= 16'h0000;
		10'h21D: instr_mem_out <= 16'h0000;
		10'h21E: instr_mem_out <= 16'h0000;
		10'h21F: instr_mem_out <= 16'h0000;
		10'h220: instr_mem_out <= 16'h0000;
		10'h221: instr_mem_out <= 16'h0000;
		10'h222: instr_mem_out <= 16'h0000;
		10'h223: instr_mem_out <= 16'h0000;
		10'h224: instr_mem_out <= 16'h0000;
		10'h225: instr_mem_out <= 16'h0000;
		10'h226: instr_mem_out <= 16'h0000;
		10'h227: instr_mem_out <= 16'h0000;
		10'h228: instr_mem_out <= 16'h0000;
		10'h229: instr_mem_out <= 16'h0000;
		10'h22A: instr_mem_out <= 16'h0000;
		10'h22B: instr_mem_out <= 16'h0000;
		10'h22C: instr_mem_out <= 16'h0000;
		10'h22D: instr_mem_out <= 16'h0000;
		10'h22E: instr_mem_out <= 16'h0000;
		10'h22F: instr_mem_out <= 16'h0000;
		10'h230: instr_mem_out <= 16'h0000;
		10'h231: instr_mem_out <= 16'h0000;
		10'h232: instr_mem_out <= 16'h0000;
		10'h233: instr_mem_out <= 16'h0000;
		10'h234: instr_mem_out <= 16'h0000;
		10'h235: instr_mem_out <= 16'h0000;
		10'h236: instr_mem_out <= 16'h0000;
		10'h237: instr_mem_out <= 16'h0000;
		10'h238: instr_mem_out <= 16'h0000;
		10'h239: instr_mem_out <= 16'h0000;
		10'h23A: instr_mem_out <= 16'h0000;
		10'h23B: instr_mem_out <= 16'h0000;
		10'h23C: instr_mem_out <= 16'h0000;
		10'h23D: instr_mem_out <= 16'h0000;
		10'h23E: instr_mem_out <= 16'h0000;
		10'h23F: instr_mem_out <= 16'h0000;
		10'h240: instr_mem_out <= 16'h0000;
		10'h241: instr_mem_out <= 16'h0000;
		10'h242: instr_mem_out <= 16'h0000;
		10'h243: instr_mem_out <= 16'h0000;
		10'h244: instr_mem_out <= 16'h0000;
		10'h245: instr_mem_out <= 16'h0000;
		10'h246: instr_mem_out <= 16'h0000;
		10'h247: instr_mem_out <= 16'h0000;
		10'h248: instr_mem_out <= 16'h0000;
		10'h249: instr_mem_out <= 16'h0000;
		10'h24A: instr_mem_out <= 16'h0000;
		10'h24B: instr_mem_out <= 16'h0000;
		10'h24C: instr_mem_out <= 16'h0000;
		10'h24D: instr_mem_out <= 16'h0000;
		10'h24E: instr_mem_out <= 16'h0000;
		10'h24F: instr_mem_out <= 16'h0000;
		10'h250: instr_mem_out <= 16'h0000;
		10'h251: instr_mem_out <= 16'h0000;
		10'h252: instr_mem_out <= 16'h0000;
		10'h253: instr_mem_out <= 16'h0000;
		10'h254: instr_mem_out <= 16'h0000;
		10'h255: instr_mem_out <= 16'h0000;
		10'h256: instr_mem_out <= 16'h0000;
		10'h257: instr_mem_out <= 16'h0000;
		10'h258: instr_mem_out <= 16'h0000;
		10'h259: instr_mem_out <= 16'h0000;
		10'h25A: instr_mem_out <= 16'h0000;
		10'h25B: instr_mem_out <= 16'h0000;
		10'h25C: instr_mem_out <= 16'h0000;
		10'h25D: instr_mem_out <= 16'h0000;
		10'h25E: instr_mem_out <= 16'h0000;
		10'h25F: instr_mem_out <= 16'h0000;
		10'h260: instr_mem_out <= 16'h0000;
		10'h261: instr_mem_out <= 16'h0000;
		10'h262: instr_mem_out <= 16'h0000;
		10'h263: instr_mem_out <= 16'h0000;
		10'h264: instr_mem_out <= 16'h0000;
		10'h265: instr_mem_out <= 16'h0000;
		10'h266: instr_mem_out <= 16'h0000;
		10'h267: instr_mem_out <= 16'h0000;
		10'h268: instr_mem_out <= 16'h0000;
		10'h269: instr_mem_out <= 16'h0000;
		10'h26A: instr_mem_out <= 16'h0000;
		10'h26B: instr_mem_out <= 16'h0000;
		10'h26C: instr_mem_out <= 16'h0000;
		10'h26D: instr_mem_out <= 16'h0000;
		10'h26E: instr_mem_out <= 16'h0000;
		10'h26F: instr_mem_out <= 16'h0000;
		10'h270: instr_mem_out <= 16'h0000;
		10'h271: instr_mem_out <= 16'h0000;
		10'h272: instr_mem_out <= 16'h0000;
		10'h273: instr_mem_out <= 16'h0000;
		10'h274: instr_mem_out <= 16'h0000;
		10'h275: instr_mem_out <= 16'h0000;
		10'h276: instr_mem_out <= 16'h0000;
		10'h277: instr_mem_out <= 16'h0000;
		10'h278: instr_mem_out <= 16'h0000;
		10'h279: instr_mem_out <= 16'h0000;
		10'h27A: instr_mem_out <= 16'h0000;
		10'h27B: instr_mem_out <= 16'h0000;
		10'h27C: instr_mem_out <= 16'h0000;
		10'h27D: instr_mem_out <= 16'h0000;
		10'h27E: instr_mem_out <= 16'h0000;
		10'h27F: instr_mem_out <= 16'h0000;
		10'h280: instr_mem_out <= 16'h0000;
		10'h281: instr_mem_out <= 16'h0000;
		10'h282: instr_mem_out <= 16'h0000;
		10'h283: instr_mem_out <= 16'h0000;
		10'h284: instr_mem_out <= 16'h0000;
		10'h285: instr_mem_out <= 16'h0000;
		10'h286: instr_mem_out <= 16'h0000;
		10'h287: instr_mem_out <= 16'h0000;
		10'h288: instr_mem_out <= 16'h0000;
		10'h289: instr_mem_out <= 16'h0000;
		10'h28A: instr_mem_out <= 16'h0000;
		10'h28B: instr_mem_out <= 16'h0000;
		10'h28C: instr_mem_out <= 16'h0000;
		10'h28D: instr_mem_out <= 16'h0000;
		10'h28E: instr_mem_out <= 16'h0000;
		10'h28F: instr_mem_out <= 16'h0000;
		10'h290: instr_mem_out <= 16'h0000;
		10'h291: instr_mem_out <= 16'h0000;
		10'h292: instr_mem_out <= 16'h0000;
		10'h293: instr_mem_out <= 16'h0000;
		10'h294: instr_mem_out <= 16'h0000;
		10'h295: instr_mem_out <= 16'h0000;
		10'h296: instr_mem_out <= 16'h0000;
		10'h297: instr_mem_out <= 16'h0000;
		10'h298: instr_mem_out <= 16'h0000;
		10'h299: instr_mem_out <= 16'h0000;
		10'h29A: instr_mem_out <= 16'h0000;
		10'h29B: instr_mem_out <= 16'h0000;
		10'h29C: instr_mem_out <= 16'h0000;
		10'h29D: instr_mem_out <= 16'h0000;
		10'h29E: instr_mem_out <= 16'h0000;
		10'h29F: instr_mem_out <= 16'h0000;
		10'h2A0: instr_mem_out <= 16'h0000;
		10'h2A1: instr_mem_out <= 16'h0000;
		10'h2A2: instr_mem_out <= 16'h0000;
		10'h2A3: instr_mem_out <= 16'h0000;
		10'h2A4: instr_mem_out <= 16'h0000;
		10'h2A5: instr_mem_out <= 16'h0000;
		10'h2A6: instr_mem_out <= 16'h0000;
		10'h2A7: instr_mem_out <= 16'h0000;
		10'h2A8: instr_mem_out <= 16'h0000;
		10'h2A9: instr_mem_out <= 16'h0000;
		10'h2AA: instr_mem_out <= 16'h0000;
		10'h2AB: instr_mem_out <= 16'h0000;
		10'h2AC: instr_mem_out <= 16'h0000;
		10'h2AD: instr_mem_out <= 16'h0000;
		10'h2AE: instr_mem_out <= 16'h0000;
		10'h2AF: instr_mem_out <= 16'h0000;
		10'h2B0: instr_mem_out <= 16'h0000;
		10'h2B1: instr_mem_out <= 16'h0000;
		10'h2B2: instr_mem_out <= 16'h0000;
		10'h2B3: instr_mem_out <= 16'h0000;
		10'h2B4: instr_mem_out <= 16'h0000;
		10'h2B5: instr_mem_out <= 16'h0000;
		10'h2B6: instr_mem_out <= 16'h0000;
		10'h2B7: instr_mem_out <= 16'h0000;
		10'h2B8: instr_mem_out <= 16'h0000;
		10'h2B9: instr_mem_out <= 16'h0000;
		10'h2BA: instr_mem_out <= 16'h0000;
		10'h2BB: instr_mem_out <= 16'h0000;
		10'h2BC: instr_mem_out <= 16'h0000;
		10'h2BD: instr_mem_out <= 16'h0000;
		10'h2BE: instr_mem_out <= 16'h0000;
		10'h2BF: instr_mem_out <= 16'h0000;
		10'h2C0: instr_mem_out <= 16'h0000;
		10'h2C1: instr_mem_out <= 16'h0000;
		10'h2C2: instr_mem_out <= 16'h0000;
		10'h2C3: instr_mem_out <= 16'h0000;
		10'h2C4: instr_mem_out <= 16'h0000;
		10'h2C5: instr_mem_out <= 16'h0000;
		10'h2C6: instr_mem_out <= 16'h0000;
		10'h2C7: instr_mem_out <= 16'h0000;
		10'h2C8: instr_mem_out <= 16'h0000;
		10'h2C9: instr_mem_out <= 16'h0000;
		10'h2CA: instr_mem_out <= 16'h0000;
		10'h2CB: instr_mem_out <= 16'h0000;
		10'h2CC: instr_mem_out <= 16'h0000;
		10'h2CD: instr_mem_out <= 16'h0000;
		10'h2CE: instr_mem_out <= 16'h0000;
		10'h2CF: instr_mem_out <= 16'h0000;
		10'h2D0: instr_mem_out <= 16'h0000;
		10'h2D1: instr_mem_out <= 16'h0000;
		10'h2D2: instr_mem_out <= 16'h0000;
		10'h2D3: instr_mem_out <= 16'h0000;
		10'h2D4: instr_mem_out <= 16'h0000;
		10'h2D5: instr_mem_out <= 16'h0000;
		10'h2D6: instr_mem_out <= 16'h0000;
		10'h2D7: instr_mem_out <= 16'h0000;
		10'h2D8: instr_mem_out <= 16'h0000;
		10'h2D9: instr_mem_out <= 16'h0000;
		10'h2DA: instr_mem_out <= 16'h0000;
		10'h2DB: instr_mem_out <= 16'h0000;
		10'h2DC: instr_mem_out <= 16'h0000;
		10'h2DD: instr_mem_out <= 16'h0000;
		10'h2DE: instr_mem_out <= 16'h0000;
		10'h2DF: instr_mem_out <= 16'h0000;
		10'h2E0: instr_mem_out <= 16'h0000;
		10'h2E1: instr_mem_out <= 16'h0000;
		10'h2E2: instr_mem_out <= 16'h0000;
		10'h2E3: instr_mem_out <= 16'h0000;
		10'h2E4: instr_mem_out <= 16'h0000;
		10'h2E5: instr_mem_out <= 16'h0000;
		10'h2E6: instr_mem_out <= 16'h0000;
		10'h2E7: instr_mem_out <= 16'h0000;
		10'h2E8: instr_mem_out <= 16'h0000;
		10'h2E9: instr_mem_out <= 16'h0000;
		10'h2EA: instr_mem_out <= 16'h0000;
		10'h2EB: instr_mem_out <= 16'h0000;
		10'h2EC: instr_mem_out <= 16'h0000;
		10'h2ED: instr_mem_out <= 16'h0000;
		10'h2EE: instr_mem_out <= 16'h0000;
		10'h2EF: instr_mem_out <= 16'h0000;
		10'h2F0: instr_mem_out <= 16'h0000;
		10'h2F1: instr_mem_out <= 16'h0000;
		10'h2F2: instr_mem_out <= 16'h0000;
		10'h2F3: instr_mem_out <= 16'h0000;
		10'h2F4: instr_mem_out <= 16'h0000;
		10'h2F5: instr_mem_out <= 16'h0000;
		10'h2F6: instr_mem_out <= 16'h0000;
		10'h2F7: instr_mem_out <= 16'h0000;
		10'h2F8: instr_mem_out <= 16'h0000;
		10'h2F9: instr_mem_out <= 16'h0000;
		10'h2FA: instr_mem_out <= 16'h0000;
		10'h2FB: instr_mem_out <= 16'h0000;
		10'h2FC: instr_mem_out <= 16'h0000;
		10'h2FD: instr_mem_out <= 16'h0000;
		10'h2FE: instr_mem_out <= 16'h0000;
		10'h2FF: instr_mem_out <= 16'h0000;
		10'h300: instr_mem_out <= 16'h0000;
		10'h301: instr_mem_out <= 16'h0000;
		10'h302: instr_mem_out <= 16'h0000;
		10'h303: instr_mem_out <= 16'h0000;
		10'h304: instr_mem_out <= 16'h0000;
		10'h305: instr_mem_out <= 16'h0000;
		10'h306: instr_mem_out <= 16'h0000;
		10'h307: instr_mem_out <= 16'h0000;
		10'h308: instr_mem_out <= 16'h0000;
		10'h309: instr_mem_out <= 16'h0000;
		10'h30A: instr_mem_out <= 16'h0000;
		10'h30B: instr_mem_out <= 16'h0000;
		10'h30C: instr_mem_out <= 16'h0000;
		10'h30D: instr_mem_out <= 16'h0000;
		10'h30E: instr_mem_out <= 16'h0000;
		10'h30F: instr_mem_out <= 16'h0000;
		10'h310: instr_mem_out <= 16'h0000;
		10'h311: instr_mem_out <= 16'h0000;
		10'h312: instr_mem_out <= 16'h0000;
		10'h313: instr_mem_out <= 16'h0000;
		10'h314: instr_mem_out <= 16'h0000;
		10'h315: instr_mem_out <= 16'h0000;
		10'h316: instr_mem_out <= 16'h0000;
		10'h317: instr_mem_out <= 16'h0000;
		10'h318: instr_mem_out <= 16'h0000;
		10'h319: instr_mem_out <= 16'h0000;
		10'h31A: instr_mem_out <= 16'h0000;
		10'h31B: instr_mem_out <= 16'h0000;
		10'h31C: instr_mem_out <= 16'h0000;
		10'h31D: instr_mem_out <= 16'h0000;
		10'h31E: instr_mem_out <= 16'h0000;
		10'h31F: instr_mem_out <= 16'h0000;
		10'h320: instr_mem_out <= 16'h0000;
		10'h321: instr_mem_out <= 16'h0000;
		10'h322: instr_mem_out <= 16'h0000;
		10'h323: instr_mem_out <= 16'h0000;
		10'h324: instr_mem_out <= 16'h0000;
		10'h325: instr_mem_out <= 16'h0000;
		10'h326: instr_mem_out <= 16'h0000;
		10'h327: instr_mem_out <= 16'h0000;
		10'h328: instr_mem_out <= 16'h0000;
		10'h329: instr_mem_out <= 16'h0000;
		10'h32A: instr_mem_out <= 16'h0000;
		10'h32B: instr_mem_out <= 16'h0000;
		10'h32C: instr_mem_out <= 16'h0000;
		10'h32D: instr_mem_out <= 16'h0000;
		10'h32E: instr_mem_out <= 16'h0000;
		10'h32F: instr_mem_out <= 16'h0000;
		10'h330: instr_mem_out <= 16'h0000;
		10'h331: instr_mem_out <= 16'h0000;
		10'h332: instr_mem_out <= 16'h0000;
		10'h333: instr_mem_out <= 16'h0000;
		10'h334: instr_mem_out <= 16'h0000;
		10'h335: instr_mem_out <= 16'h0000;
		10'h336: instr_mem_out <= 16'h0000;
		10'h337: instr_mem_out <= 16'h0000;
		10'h338: instr_mem_out <= 16'h0000;
		10'h339: instr_mem_out <= 16'h0000;
		10'h33A: instr_mem_out <= 16'h0000;
		10'h33B: instr_mem_out <= 16'h0000;
		10'h33C: instr_mem_out <= 16'h0000;
		10'h33D: instr_mem_out <= 16'h0000;
		10'h33E: instr_mem_out <= 16'h0000;
		10'h33F: instr_mem_out <= 16'h0000;
		10'h340: instr_mem_out <= 16'h0000;
		10'h341: instr_mem_out <= 16'h0000;
		10'h342: instr_mem_out <= 16'h0000;
		10'h343: instr_mem_out <= 16'h0000;
		10'h344: instr_mem_out <= 16'h0000;
		10'h345: instr_mem_out <= 16'h0000;
		10'h346: instr_mem_out <= 16'h0000;
		10'h347: instr_mem_out <= 16'h0000;
		10'h348: instr_mem_out <= 16'h0000;
		10'h349: instr_mem_out <= 16'h0000;
		10'h34A: instr_mem_out <= 16'h0000;
		10'h34B: instr_mem_out <= 16'h0000;
		10'h34C: instr_mem_out <= 16'h0000;
		10'h34D: instr_mem_out <= 16'h0000;
		10'h34E: instr_mem_out <= 16'h0000;
		10'h34F: instr_mem_out <= 16'h0000;
		10'h350: instr_mem_out <= 16'h0000;
		10'h351: instr_mem_out <= 16'h0000;
		10'h352: instr_mem_out <= 16'h0000;
		10'h353: instr_mem_out <= 16'h0000;
		10'h354: instr_mem_out <= 16'h0000;
		10'h355: instr_mem_out <= 16'h0000;
		10'h356: instr_mem_out <= 16'h0000;
		10'h357: instr_mem_out <= 16'h0000;
		10'h358: instr_mem_out <= 16'h0000;
		10'h359: instr_mem_out <= 16'h0000;
		10'h35A: instr_mem_out <= 16'h0000;
		10'h35B: instr_mem_out <= 16'h0000;
		10'h35C: instr_mem_out <= 16'h0000;
		10'h35D: instr_mem_out <= 16'h0000;
		10'h35E: instr_mem_out <= 16'h0000;
		10'h35F: instr_mem_out <= 16'h0000;
		10'h360: instr_mem_out <= 16'h0000;
		10'h361: instr_mem_out <= 16'h0000;
		10'h362: instr_mem_out <= 16'h0000;
		10'h363: instr_mem_out <= 16'h0000;
		10'h364: instr_mem_out <= 16'h0000;
		10'h365: instr_mem_out <= 16'h0000;
		10'h366: instr_mem_out <= 16'h0000;
		10'h367: instr_mem_out <= 16'h0000;
		10'h368: instr_mem_out <= 16'h0000;
		10'h369: instr_mem_out <= 16'h0000;
		10'h36A: instr_mem_out <= 16'h0000;
		10'h36B: instr_mem_out <= 16'h0000;
		10'h36C: instr_mem_out <= 16'h0000;
		10'h36D: instr_mem_out <= 16'h0000;
		10'h36E: instr_mem_out <= 16'h0000;
		10'h36F: instr_mem_out <= 16'h0000;
		10'h370: instr_mem_out <= 16'h0000;
		10'h371: instr_mem_out <= 16'h0000;
		10'h372: instr_mem_out <= 16'h0000;
		10'h373: instr_mem_out <= 16'h0000;
		10'h374: instr_mem_out <= 16'h0000;
		10'h375: instr_mem_out <= 16'h0000;
		10'h376: instr_mem_out <= 16'h0000;
		10'h377: instr_mem_out <= 16'h0000;
		10'h378: instr_mem_out <= 16'h0000;
		10'h379: instr_mem_out <= 16'h0000;
		10'h37A: instr_mem_out <= 16'h0000;
		10'h37B: instr_mem_out <= 16'h0000;
		10'h37C: instr_mem_out <= 16'h0000;
		10'h37D: instr_mem_out <= 16'h0000;
		10'h37E: instr_mem_out <= 16'h0000;
		10'h37F: instr_mem_out <= 16'h0000;
		10'h380: instr_mem_out <= 16'h0000;
		10'h381: instr_mem_out <= 16'h0000;
		10'h382: instr_mem_out <= 16'h0000;
		10'h383: instr_mem_out <= 16'h0000;
		10'h384: instr_mem_out <= 16'h0000;
		10'h385: instr_mem_out <= 16'h0000;
		10'h386: instr_mem_out <= 16'h0000;
		10'h387: instr_mem_out <= 16'h0000;
		10'h388: instr_mem_out <= 16'h0000;
		10'h389: instr_mem_out <= 16'h0000;
		10'h38A: instr_mem_out <= 16'h0000;
		10'h38B: instr_mem_out <= 16'h0000;
		10'h38C: instr_mem_out <= 16'h0000;
		10'h38D: instr_mem_out <= 16'h0000;
		10'h38E: instr_mem_out <= 16'h0000;
		10'h38F: instr_mem_out <= 16'h0000;
		10'h390: instr_mem_out <= 16'h0000;
		10'h391: instr_mem_out <= 16'h0000;
		10'h392: instr_mem_out <= 16'h0000;
		10'h393: instr_mem_out <= 16'h0000;
		10'h394: instr_mem_out <= 16'h0000;
		10'h395: instr_mem_out <= 16'h0000;
		10'h396: instr_mem_out <= 16'h0000;
		10'h397: instr_mem_out <= 16'h0000;
		10'h398: instr_mem_out <= 16'h0000;
		10'h399: instr_mem_out <= 16'h0000;
		10'h39A: instr_mem_out <= 16'h0000;
		10'h39B: instr_mem_out <= 16'h0000;
		10'h39C: instr_mem_out <= 16'h0000;
		10'h39D: instr_mem_out <= 16'h0000;
		10'h39E: instr_mem_out <= 16'h0000;
		10'h39F: instr_mem_out <= 16'h0000;
		10'h3A0: instr_mem_out <= 16'h0000;
		10'h3A1: instr_mem_out <= 16'h0000;
		10'h3A2: instr_mem_out <= 16'h0000;
		10'h3A3: instr_mem_out <= 16'h0000;
		10'h3A4: instr_mem_out <= 16'h0000;
		10'h3A5: instr_mem_out <= 16'h0000;
		10'h3A6: instr_mem_out <= 16'h0000;
		10'h3A7: instr_mem_out <= 16'h0000;
		10'h3A8: instr_mem_out <= 16'h0000;
		10'h3A9: instr_mem_out <= 16'h0000;
		10'h3AA: instr_mem_out <= 16'h0000;
		10'h3AB: instr_mem_out <= 16'h0000;
		10'h3AC: instr_mem_out <= 16'h0000;
		10'h3AD: instr_mem_out <= 16'h0000;
		10'h3AE: instr_mem_out <= 16'h0000;
		10'h3AF: instr_mem_out <= 16'h0000;
		10'h3B0: instr_mem_out <= 16'h0000;
		10'h3B1: instr_mem_out <= 16'h0000;
		10'h3B2: instr_mem_out <= 16'h0000;
		10'h3B3: instr_mem_out <= 16'h0000;
		10'h3B4: instr_mem_out <= 16'h0000;
		10'h3B5: instr_mem_out <= 16'h0000;
		10'h3B6: instr_mem_out <= 16'h0000;
		10'h3B7: instr_mem_out <= 16'h0000;
		10'h3B8: instr_mem_out <= 16'h0000;
		10'h3B9: instr_mem_out <= 16'h0000;
		10'h3BA: instr_mem_out <= 16'h0000;
		10'h3BB: instr_mem_out <= 16'h0000;
		10'h3BC: instr_mem_out <= 16'h0000;
		10'h3BD: instr_mem_out <= 16'h0000;
		10'h3BE: instr_mem_out <= 16'h0000;
		10'h3BF: instr_mem_out <= 16'h0000;
		10'h3C0: instr_mem_out <= 16'h0000;
		10'h3C1: instr_mem_out <= 16'h0000;
		10'h3C2: instr_mem_out <= 16'h0000;
		10'h3C3: instr_mem_out <= 16'h0000;
		10'h3C4: instr_mem_out <= 16'h0000;
		10'h3C5: instr_mem_out <= 16'h0000;
		10'h3C6: instr_mem_out <= 16'h0000;
		10'h3C7: instr_mem_out <= 16'h0000;
		10'h3C8: instr_mem_out <= 16'h0000;
		10'h3C9: instr_mem_out <= 16'h0000;
		10'h3CA: instr_mem_out <= 16'h0000;
		10'h3CB: instr_mem_out <= 16'h0000;
		10'h3CC: instr_mem_out <= 16'h0000;
		10'h3CD: instr_mem_out <= 16'h0000;
		10'h3CE: instr_mem_out <= 16'h0000;
		10'h3CF: instr_mem_out <= 16'h0000;
		10'h3D0: instr_mem_out <= 16'h0000;
		10'h3D1: instr_mem_out <= 16'h0000;
		10'h3D2: instr_mem_out <= 16'h0000;
		10'h3D3: instr_mem_out <= 16'h0000;
		10'h3D4: instr_mem_out <= 16'h0000;
		10'h3D5: instr_mem_out <= 16'h0000;
		10'h3D6: instr_mem_out <= 16'h0000;
		10'h3D7: instr_mem_out <= 16'h0000;
		10'h3D8: instr_mem_out <= 16'h0000;
		10'h3D9: instr_mem_out <= 16'h0000;
		10'h3DA: instr_mem_out <= 16'h0000;
		10'h3DB: instr_mem_out <= 16'h0000;
		10'h3DC: instr_mem_out <= 16'h0000;
		10'h3DD: instr_mem_out <= 16'h0000;
		10'h3DE: instr_mem_out <= 16'h0000;
		10'h3DF: instr_mem_out <= 16'h0000;
		10'h3E0: instr_mem_out <= 16'h0000;
		10'h3E1: instr_mem_out <= 16'h0000;
		10'h3E2: instr_mem_out <= 16'h0000;
		10'h3E3: instr_mem_out <= 16'h0000;
		10'h3E4: instr_mem_out <= 16'h0000;
		10'h3E5: instr_mem_out <= 16'h0000;
		10'h3E6: instr_mem_out <= 16'h0000;
		10'h3E7: instr_mem_out <= 16'h0000;
		10'h3E8: instr_mem_out <= 16'h0000;
		10'h3E9: instr_mem_out <= 16'h0000;
		10'h3EA: instr_mem_out <= 16'h0000;
		10'h3EB: instr_mem_out <= 16'h0000;
		10'h3EC: instr_mem_out <= 16'h0000;
		10'h3ED: instr_mem_out <= 16'h0000;
		10'h3EE: instr_mem_out <= 16'h0000;
		10'h3EF: instr_mem_out <= 16'h0000;
		10'h3F0: instr_mem_out <= 16'h0000;
		10'h3F1: instr_mem_out <= 16'h0000;
		10'h3F2: instr_mem_out <= 16'h0000;
		10'h3F3: instr_mem_out <= 16'h0000;
		10'h3F4: instr_mem_out <= 16'h0000;
		10'h3F5: instr_mem_out <= 16'h0000;
		10'h3F6: instr_mem_out <= 16'h0000;
		10'h3F7: instr_mem_out <= 16'h0000;
		10'h3F8: instr_mem_out <= 16'h0000;
		10'h3F9: instr_mem_out <= 16'h0000;
		10'h3FA: instr_mem_out <= 16'h0000;
		10'h3FB: instr_mem_out <= 16'h0000;
		10'h3FC: instr_mem_out <= 16'h0000;
		10'h3FD: instr_mem_out <= 16'h0000;
		10'h3FE: instr_mem_out <= 16'h0000;
		10'h3FF: instr_mem_out <= 16'h0000;
		default: instr_mem_out <= 16'h0000;
	endcase
end
endmodule
