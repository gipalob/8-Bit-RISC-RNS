module Instr_Mem #(parameter PROG_CTR_WID = 10) (
	input [PROG_CTR_WID-1:0] prog_ctr,
	output reg [15:0] instruction
);
always @(*) begin
	case (prog_ctr)
		10'h000: instruction <= 16'h9008;
		10'h001: instruction <= 16'h9102;
		10'h002: instruction <= 16'hA810;
		10'h003: instruction <= 16'h0000;
		10'h004: instruction <= 16'h9910;
		10'h005: instruction <= 16'h0000;
		10'h006: instruction <= 16'hA210;
		10'h007: instruction <= 16'h0000;
		10'h008: instruction <= 16'h920A;
		10'h009: instruction <= 16'hAB28;
		10'h00A: instruction <= 16'hACAB;
		10'h00B: instruction <= 16'h0000;
		10'h00C: instruction <= 16'hBB0C;
		10'h00D: instruction <= 16'hC40C;
		10'h00E: instruction <= 16'hCD10;
		10'h00F: instruction <= 16'h0000;
		10'h010: instruction <= 16'h0000;
		10'h011: instruction <= 16'h0000;
		10'h012: instruction <= 16'h0000;
		10'h013: instruction <= 16'h0000;
		10'h014: instruction <= 16'h0000;
		10'h015: instruction <= 16'h0000;
		10'h016: instruction <= 16'h0000;
		10'h017: instruction <= 16'h0000;
		10'h018: instruction <= 16'h0000;
		10'h019: instruction <= 16'h0000;
		10'h01A: instruction <= 16'h0000;
		10'h01B: instruction <= 16'h0000;
		10'h01C: instruction <= 16'h0000;
		10'h01D: instruction <= 16'h0000;
		10'h01E: instruction <= 16'h0000;
		10'h01F: instruction <= 16'h0000;
		10'h020: instruction <= 16'h0000;
		10'h021: instruction <= 16'h0000;
		10'h022: instruction <= 16'h0000;
		10'h023: instruction <= 16'h0000;
		10'h024: instruction <= 16'h0000;
		10'h025: instruction <= 16'h0000;
		10'h026: instruction <= 16'h0000;
		10'h027: instruction <= 16'h0000;
		10'h028: instruction <= 16'h0000;
		10'h029: instruction <= 16'h0000;
		10'h02A: instruction <= 16'h0000;
		10'h02B: instruction <= 16'h0000;
		10'h02C: instruction <= 16'h0000;
		10'h02D: instruction <= 16'h0000;
		10'h02E: instruction <= 16'h0000;
		10'h02F: instruction <= 16'h0000;
		10'h030: instruction <= 16'h0000;
		10'h031: instruction <= 16'h0000;
		10'h032: instruction <= 16'h0000;
		10'h033: instruction <= 16'h0000;
		10'h034: instruction <= 16'h0000;
		10'h035: instruction <= 16'h0000;
		10'h036: instruction <= 16'h0000;
		10'h037: instruction <= 16'h0000;
		10'h038: instruction <= 16'h0000;
		10'h039: instruction <= 16'h0000;
		10'h03A: instruction <= 16'h0000;
		10'h03B: instruction <= 16'h0000;
		10'h03C: instruction <= 16'h0000;
		10'h03D: instruction <= 16'h0000;
		10'h03E: instruction <= 16'h0000;
		10'h03F: instruction <= 16'h0000;
		10'h040: instruction <= 16'h0000;
		10'h041: instruction <= 16'h0000;
		10'h042: instruction <= 16'h0000;
		10'h043: instruction <= 16'h0000;
		10'h044: instruction <= 16'h0000;
		10'h045: instruction <= 16'h0000;
		10'h046: instruction <= 16'h0000;
		10'h047: instruction <= 16'h0000;
		10'h048: instruction <= 16'h0000;
		10'h049: instruction <= 16'h0000;
		10'h04A: instruction <= 16'h0000;
		10'h04B: instruction <= 16'h0000;
		10'h04C: instruction <= 16'h0000;
		10'h04D: instruction <= 16'h0000;
		10'h04E: instruction <= 16'h0000;
		10'h04F: instruction <= 16'h0000;
		10'h050: instruction <= 16'h0000;
		10'h051: instruction <= 16'h0000;
		10'h052: instruction <= 16'h0000;
		10'h053: instruction <= 16'h0000;
		10'h054: instruction <= 16'h0000;
		10'h055: instruction <= 16'h0000;
		10'h056: instruction <= 16'h0000;
		10'h057: instruction <= 16'h0000;
		10'h058: instruction <= 16'h0000;
		10'h059: instruction <= 16'h0000;
		10'h05A: instruction <= 16'h0000;
		10'h05B: instruction <= 16'h0000;
		10'h05C: instruction <= 16'h0000;
		10'h05D: instruction <= 16'h0000;
		10'h05E: instruction <= 16'h0000;
		10'h05F: instruction <= 16'h0000;
		10'h060: instruction <= 16'h0000;
		10'h061: instruction <= 16'h0000;
		10'h062: instruction <= 16'h0000;
		10'h063: instruction <= 16'h0000;
		10'h064: instruction <= 16'h0000;
		10'h065: instruction <= 16'h0000;
		10'h066: instruction <= 16'h0000;
		10'h067: instruction <= 16'h0000;
		10'h068: instruction <= 16'h0000;
		10'h069: instruction <= 16'h0000;
		10'h06A: instruction <= 16'h0000;
		10'h06B: instruction <= 16'h0000;
		10'h06C: instruction <= 16'h0000;
		10'h06D: instruction <= 16'h0000;
		10'h06E: instruction <= 16'h0000;
		10'h06F: instruction <= 16'h0000;
		10'h070: instruction <= 16'h0000;
		10'h071: instruction <= 16'h0000;
		10'h072: instruction <= 16'h0000;
		10'h073: instruction <= 16'h0000;
		10'h074: instruction <= 16'h0000;
		10'h075: instruction <= 16'h0000;
		10'h076: instruction <= 16'h0000;
		10'h077: instruction <= 16'h0000;
		10'h078: instruction <= 16'h0000;
		10'h079: instruction <= 16'h0000;
		10'h07A: instruction <= 16'h0000;
		10'h07B: instruction <= 16'h0000;
		10'h07C: instruction <= 16'h0000;
		10'h07D: instruction <= 16'h0000;
		10'h07E: instruction <= 16'h0000;
		10'h07F: instruction <= 16'h0000;
		10'h080: instruction <= 16'h0000;
		10'h081: instruction <= 16'h0000;
		10'h082: instruction <= 16'h0000;
		10'h083: instruction <= 16'h0000;
		10'h084: instruction <= 16'h0000;
		10'h085: instruction <= 16'h0000;
		10'h086: instruction <= 16'h0000;
		10'h087: instruction <= 16'h0000;
		10'h088: instruction <= 16'h0000;
		10'h089: instruction <= 16'h0000;
		10'h08A: instruction <= 16'h0000;
		10'h08B: instruction <= 16'h0000;
		10'h08C: instruction <= 16'h0000;
		10'h08D: instruction <= 16'h0000;
		10'h08E: instruction <= 16'h0000;
		10'h08F: instruction <= 16'h0000;
		10'h090: instruction <= 16'h0000;
		10'h091: instruction <= 16'h0000;
		10'h092: instruction <= 16'h0000;
		10'h093: instruction <= 16'h0000;
		10'h094: instruction <= 16'h0000;
		10'h095: instruction <= 16'h0000;
		10'h096: instruction <= 16'h0000;
		10'h097: instruction <= 16'h0000;
		10'h098: instruction <= 16'h0000;
		10'h099: instruction <= 16'h0000;
		10'h09A: instruction <= 16'h0000;
		10'h09B: instruction <= 16'h0000;
		10'h09C: instruction <= 16'h0000;
		10'h09D: instruction <= 16'h0000;
		10'h09E: instruction <= 16'h0000;
		10'h09F: instruction <= 16'h0000;
		10'h0A0: instruction <= 16'h0000;
		10'h0A1: instruction <= 16'h0000;
		10'h0A2: instruction <= 16'h0000;
		10'h0A3: instruction <= 16'h0000;
		10'h0A4: instruction <= 16'h0000;
		10'h0A5: instruction <= 16'h0000;
		10'h0A6: instruction <= 16'h0000;
		10'h0A7: instruction <= 16'h0000;
		10'h0A8: instruction <= 16'h0000;
		10'h0A9: instruction <= 16'h0000;
		10'h0AA: instruction <= 16'h0000;
		10'h0AB: instruction <= 16'h0000;
		10'h0AC: instruction <= 16'h0000;
		10'h0AD: instruction <= 16'h0000;
		10'h0AE: instruction <= 16'h0000;
		10'h0AF: instruction <= 16'h0000;
		10'h0B0: instruction <= 16'h0000;
		10'h0B1: instruction <= 16'h0000;
		10'h0B2: instruction <= 16'h0000;
		10'h0B3: instruction <= 16'h0000;
		10'h0B4: instruction <= 16'h0000;
		10'h0B5: instruction <= 16'h0000;
		10'h0B6: instruction <= 16'h0000;
		10'h0B7: instruction <= 16'h0000;
		10'h0B8: instruction <= 16'h0000;
		10'h0B9: instruction <= 16'h0000;
		10'h0BA: instruction <= 16'h0000;
		10'h0BB: instruction <= 16'h0000;
		10'h0BC: instruction <= 16'h0000;
		10'h0BD: instruction <= 16'h0000;
		10'h0BE: instruction <= 16'h0000;
		10'h0BF: instruction <= 16'h0000;
		10'h0C0: instruction <= 16'h0000;
		10'h0C1: instruction <= 16'h0000;
		10'h0C2: instruction <= 16'h0000;
		10'h0C3: instruction <= 16'h0000;
		10'h0C4: instruction <= 16'h0000;
		10'h0C5: instruction <= 16'h0000;
		10'h0C6: instruction <= 16'h0000;
		10'h0C7: instruction <= 16'h0000;
		10'h0C8: instruction <= 16'h0000;
		10'h0C9: instruction <= 16'h0000;
		10'h0CA: instruction <= 16'h0000;
		10'h0CB: instruction <= 16'h0000;
		10'h0CC: instruction <= 16'h0000;
		10'h0CD: instruction <= 16'h0000;
		10'h0CE: instruction <= 16'h0000;
		10'h0CF: instruction <= 16'h0000;
		10'h0D0: instruction <= 16'h0000;
		10'h0D1: instruction <= 16'h0000;
		10'h0D2: instruction <= 16'h0000;
		10'h0D3: instruction <= 16'h0000;
		10'h0D4: instruction <= 16'h0000;
		10'h0D5: instruction <= 16'h0000;
		10'h0D6: instruction <= 16'h0000;
		10'h0D7: instruction <= 16'h0000;
		10'h0D8: instruction <= 16'h0000;
		10'h0D9: instruction <= 16'h0000;
		10'h0DA: instruction <= 16'h0000;
		10'h0DB: instruction <= 16'h0000;
		10'h0DC: instruction <= 16'h0000;
		10'h0DD: instruction <= 16'h0000;
		10'h0DE: instruction <= 16'h0000;
		10'h0DF: instruction <= 16'h0000;
		10'h0E0: instruction <= 16'h0000;
		10'h0E1: instruction <= 16'h0000;
		10'h0E2: instruction <= 16'h0000;
		10'h0E3: instruction <= 16'h0000;
		10'h0E4: instruction <= 16'h0000;
		10'h0E5: instruction <= 16'h0000;
		10'h0E6: instruction <= 16'h0000;
		10'h0E7: instruction <= 16'h0000;
		10'h0E8: instruction <= 16'h0000;
		10'h0E9: instruction <= 16'h0000;
		10'h0EA: instruction <= 16'h0000;
		10'h0EB: instruction <= 16'h0000;
		10'h0EC: instruction <= 16'h0000;
		10'h0ED: instruction <= 16'h0000;
		10'h0EE: instruction <= 16'h0000;
		10'h0EF: instruction <= 16'h0000;
		10'h0F0: instruction <= 16'h0000;
		10'h0F1: instruction <= 16'h0000;
		10'h0F2: instruction <= 16'h0000;
		10'h0F3: instruction <= 16'h0000;
		10'h0F4: instruction <= 16'h0000;
		10'h0F5: instruction <= 16'h0000;
		10'h0F6: instruction <= 16'h0000;
		10'h0F7: instruction <= 16'h0000;
		10'h0F8: instruction <= 16'h0000;
		10'h0F9: instruction <= 16'h0000;
		10'h0FA: instruction <= 16'h0000;
		10'h0FB: instruction <= 16'h0000;
		10'h0FC: instruction <= 16'h0000;
		10'h0FD: instruction <= 16'h0000;
		10'h0FE: instruction <= 16'h0000;
		10'h0FF: instruction <= 16'h0000;
		10'h100: instruction <= 16'h0000;
		10'h101: instruction <= 16'h0000;
		10'h102: instruction <= 16'h0000;
		10'h103: instruction <= 16'h0000;
		10'h104: instruction <= 16'h0000;
		10'h105: instruction <= 16'h0000;
		10'h106: instruction <= 16'h0000;
		10'h107: instruction <= 16'h0000;
		10'h108: instruction <= 16'h0000;
		10'h109: instruction <= 16'h0000;
		10'h10A: instruction <= 16'h0000;
		10'h10B: instruction <= 16'h0000;
		10'h10C: instruction <= 16'h0000;
		10'h10D: instruction <= 16'h0000;
		10'h10E: instruction <= 16'h0000;
		10'h10F: instruction <= 16'h0000;
		10'h110: instruction <= 16'h0000;
		10'h111: instruction <= 16'h0000;
		10'h112: instruction <= 16'h0000;
		10'h113: instruction <= 16'h0000;
		10'h114: instruction <= 16'h0000;
		10'h115: instruction <= 16'h0000;
		10'h116: instruction <= 16'h0000;
		10'h117: instruction <= 16'h0000;
		10'h118: instruction <= 16'h0000;
		10'h119: instruction <= 16'h0000;
		10'h11A: instruction <= 16'h0000;
		10'h11B: instruction <= 16'h0000;
		10'h11C: instruction <= 16'h0000;
		10'h11D: instruction <= 16'h0000;
		10'h11E: instruction <= 16'h0000;
		10'h11F: instruction <= 16'h0000;
		10'h120: instruction <= 16'h0000;
		10'h121: instruction <= 16'h0000;
		10'h122: instruction <= 16'h0000;
		10'h123: instruction <= 16'h0000;
		10'h124: instruction <= 16'h0000;
		10'h125: instruction <= 16'h0000;
		10'h126: instruction <= 16'h0000;
		10'h127: instruction <= 16'h0000;
		10'h128: instruction <= 16'h0000;
		10'h129: instruction <= 16'h0000;
		10'h12A: instruction <= 16'h0000;
		10'h12B: instruction <= 16'h0000;
		10'h12C: instruction <= 16'h0000;
		10'h12D: instruction <= 16'h0000;
		10'h12E: instruction <= 16'h0000;
		10'h12F: instruction <= 16'h0000;
		10'h130: instruction <= 16'h0000;
		10'h131: instruction <= 16'h0000;
		10'h132: instruction <= 16'h0000;
		10'h133: instruction <= 16'h0000;
		10'h134: instruction <= 16'h0000;
		10'h135: instruction <= 16'h0000;
		10'h136: instruction <= 16'h0000;
		10'h137: instruction <= 16'h0000;
		10'h138: instruction <= 16'h0000;
		10'h139: instruction <= 16'h0000;
		10'h13A: instruction <= 16'h0000;
		10'h13B: instruction <= 16'h0000;
		10'h13C: instruction <= 16'h0000;
		10'h13D: instruction <= 16'h0000;
		10'h13E: instruction <= 16'h0000;
		10'h13F: instruction <= 16'h0000;
		10'h140: instruction <= 16'h0000;
		10'h141: instruction <= 16'h0000;
		10'h142: instruction <= 16'h0000;
		10'h143: instruction <= 16'h0000;
		10'h144: instruction <= 16'h0000;
		10'h145: instruction <= 16'h0000;
		10'h146: instruction <= 16'h0000;
		10'h147: instruction <= 16'h0000;
		10'h148: instruction <= 16'h0000;
		10'h149: instruction <= 16'h0000;
		10'h14A: instruction <= 16'h0000;
		10'h14B: instruction <= 16'h0000;
		10'h14C: instruction <= 16'h0000;
		10'h14D: instruction <= 16'h0000;
		10'h14E: instruction <= 16'h0000;
		10'h14F: instruction <= 16'h0000;
		10'h150: instruction <= 16'h0000;
		10'h151: instruction <= 16'h0000;
		10'h152: instruction <= 16'h0000;
		10'h153: instruction <= 16'h0000;
		10'h154: instruction <= 16'h0000;
		10'h155: instruction <= 16'h0000;
		10'h156: instruction <= 16'h0000;
		10'h157: instruction <= 16'h0000;
		10'h158: instruction <= 16'h0000;
		10'h159: instruction <= 16'h0000;
		10'h15A: instruction <= 16'h0000;
		10'h15B: instruction <= 16'h0000;
		10'h15C: instruction <= 16'h0000;
		10'h15D: instruction <= 16'h0000;
		10'h15E: instruction <= 16'h0000;
		10'h15F: instruction <= 16'h0000;
		10'h160: instruction <= 16'h0000;
		10'h161: instruction <= 16'h0000;
		10'h162: instruction <= 16'h0000;
		10'h163: instruction <= 16'h0000;
		10'h164: instruction <= 16'h0000;
		10'h165: instruction <= 16'h0000;
		10'h166: instruction <= 16'h0000;
		10'h167: instruction <= 16'h0000;
		10'h168: instruction <= 16'h0000;
		10'h169: instruction <= 16'h0000;
		10'h16A: instruction <= 16'h0000;
		10'h16B: instruction <= 16'h0000;
		10'h16C: instruction <= 16'h0000;
		10'h16D: instruction <= 16'h0000;
		10'h16E: instruction <= 16'h0000;
		10'h16F: instruction <= 16'h0000;
		10'h170: instruction <= 16'h0000;
		10'h171: instruction <= 16'h0000;
		10'h172: instruction <= 16'h0000;
		10'h173: instruction <= 16'h0000;
		10'h174: instruction <= 16'h0000;
		10'h175: instruction <= 16'h0000;
		10'h176: instruction <= 16'h0000;
		10'h177: instruction <= 16'h0000;
		10'h178: instruction <= 16'h0000;
		10'h179: instruction <= 16'h0000;
		10'h17A: instruction <= 16'h0000;
		10'h17B: instruction <= 16'h0000;
		10'h17C: instruction <= 16'h0000;
		10'h17D: instruction <= 16'h0000;
		10'h17E: instruction <= 16'h0000;
		10'h17F: instruction <= 16'h0000;
		10'h180: instruction <= 16'h0000;
		10'h181: instruction <= 16'h0000;
		10'h182: instruction <= 16'h0000;
		10'h183: instruction <= 16'h0000;
		10'h184: instruction <= 16'h0000;
		10'h185: instruction <= 16'h0000;
		10'h186: instruction <= 16'h0000;
		10'h187: instruction <= 16'h0000;
		10'h188: instruction <= 16'h0000;
		10'h189: instruction <= 16'h0000;
		10'h18A: instruction <= 16'h0000;
		10'h18B: instruction <= 16'h0000;
		10'h18C: instruction <= 16'h0000;
		10'h18D: instruction <= 16'h0000;
		10'h18E: instruction <= 16'h0000;
		10'h18F: instruction <= 16'h0000;
		10'h190: instruction <= 16'h0000;
		10'h191: instruction <= 16'h0000;
		10'h192: instruction <= 16'h0000;
		10'h193: instruction <= 16'h0000;
		10'h194: instruction <= 16'h0000;
		10'h195: instruction <= 16'h0000;
		10'h196: instruction <= 16'h0000;
		10'h197: instruction <= 16'h0000;
		10'h198: instruction <= 16'h0000;
		10'h199: instruction <= 16'h0000;
		10'h19A: instruction <= 16'h0000;
		10'h19B: instruction <= 16'h0000;
		10'h19C: instruction <= 16'h0000;
		10'h19D: instruction <= 16'h0000;
		10'h19E: instruction <= 16'h0000;
		10'h19F: instruction <= 16'h0000;
		10'h1A0: instruction <= 16'h0000;
		10'h1A1: instruction <= 16'h0000;
		10'h1A2: instruction <= 16'h0000;
		10'h1A3: instruction <= 16'h0000;
		10'h1A4: instruction <= 16'h0000;
		10'h1A5: instruction <= 16'h0000;
		10'h1A6: instruction <= 16'h0000;
		10'h1A7: instruction <= 16'h0000;
		10'h1A8: instruction <= 16'h0000;
		10'h1A9: instruction <= 16'h0000;
		10'h1AA: instruction <= 16'h0000;
		10'h1AB: instruction <= 16'h0000;
		10'h1AC: instruction <= 16'h0000;
		10'h1AD: instruction <= 16'h0000;
		10'h1AE: instruction <= 16'h0000;
		10'h1AF: instruction <= 16'h0000;
		10'h1B0: instruction <= 16'h0000;
		10'h1B1: instruction <= 16'h0000;
		10'h1B2: instruction <= 16'h0000;
		10'h1B3: instruction <= 16'h0000;
		10'h1B4: instruction <= 16'h0000;
		10'h1B5: instruction <= 16'h0000;
		10'h1B6: instruction <= 16'h0000;
		10'h1B7: instruction <= 16'h0000;
		10'h1B8: instruction <= 16'h0000;
		10'h1B9: instruction <= 16'h0000;
		10'h1BA: instruction <= 16'h0000;
		10'h1BB: instruction <= 16'h0000;
		10'h1BC: instruction <= 16'h0000;
		10'h1BD: instruction <= 16'h0000;
		10'h1BE: instruction <= 16'h0000;
		10'h1BF: instruction <= 16'h0000;
		10'h1C0: instruction <= 16'h0000;
		10'h1C1: instruction <= 16'h0000;
		10'h1C2: instruction <= 16'h0000;
		10'h1C3: instruction <= 16'h0000;
		10'h1C4: instruction <= 16'h0000;
		10'h1C5: instruction <= 16'h0000;
		10'h1C6: instruction <= 16'h0000;
		10'h1C7: instruction <= 16'h0000;
		10'h1C8: instruction <= 16'h0000;
		10'h1C9: instruction <= 16'h0000;
		10'h1CA: instruction <= 16'h0000;
		10'h1CB: instruction <= 16'h0000;
		10'h1CC: instruction <= 16'h0000;
		10'h1CD: instruction <= 16'h0000;
		10'h1CE: instruction <= 16'h0000;
		10'h1CF: instruction <= 16'h0000;
		10'h1D0: instruction <= 16'h0000;
		10'h1D1: instruction <= 16'h0000;
		10'h1D2: instruction <= 16'h0000;
		10'h1D3: instruction <= 16'h0000;
		10'h1D4: instruction <= 16'h0000;
		10'h1D5: instruction <= 16'h0000;
		10'h1D6: instruction <= 16'h0000;
		10'h1D7: instruction <= 16'h0000;
		10'h1D8: instruction <= 16'h0000;
		10'h1D9: instruction <= 16'h0000;
		10'h1DA: instruction <= 16'h0000;
		10'h1DB: instruction <= 16'h0000;
		10'h1DC: instruction <= 16'h0000;
		10'h1DD: instruction <= 16'h0000;
		10'h1DE: instruction <= 16'h0000;
		10'h1DF: instruction <= 16'h0000;
		10'h1E0: instruction <= 16'h0000;
		10'h1E1: instruction <= 16'h0000;
		10'h1E2: instruction <= 16'h0000;
		10'h1E3: instruction <= 16'h0000;
		10'h1E4: instruction <= 16'h0000;
		10'h1E5: instruction <= 16'h0000;
		10'h1E6: instruction <= 16'h0000;
		10'h1E7: instruction <= 16'h0000;
		10'h1E8: instruction <= 16'h0000;
		10'h1E9: instruction <= 16'h0000;
		10'h1EA: instruction <= 16'h0000;
		10'h1EB: instruction <= 16'h0000;
		10'h1EC: instruction <= 16'h0000;
		10'h1ED: instruction <= 16'h0000;
		10'h1EE: instruction <= 16'h0000;
		10'h1EF: instruction <= 16'h0000;
		10'h1F0: instruction <= 16'h0000;
		10'h1F1: instruction <= 16'h0000;
		10'h1F2: instruction <= 16'h0000;
		10'h1F3: instruction <= 16'h0000;
		10'h1F4: instruction <= 16'h0000;
		10'h1F5: instruction <= 16'h0000;
		10'h1F6: instruction <= 16'h0000;
		10'h1F7: instruction <= 16'h0000;
		10'h1F8: instruction <= 16'h0000;
		10'h1F9: instruction <= 16'h0000;
		10'h1FA: instruction <= 16'h0000;
		10'h1FB: instruction <= 16'h0000;
		10'h1FC: instruction <= 16'h0000;
		10'h1FD: instruction <= 16'h0000;
		10'h1FE: instruction <= 16'h0000;
		10'h1FF: instruction <= 16'h0000;
		10'h200: instruction <= 16'h0000;
		10'h201: instruction <= 16'h0000;
		10'h202: instruction <= 16'h0000;
		10'h203: instruction <= 16'h0000;
		10'h204: instruction <= 16'h0000;
		10'h205: instruction <= 16'h0000;
		10'h206: instruction <= 16'h0000;
		10'h207: instruction <= 16'h0000;
		10'h208: instruction <= 16'h0000;
		10'h209: instruction <= 16'h0000;
		10'h20A: instruction <= 16'h0000;
		10'h20B: instruction <= 16'h0000;
		10'h20C: instruction <= 16'h0000;
		10'h20D: instruction <= 16'h0000;
		10'h20E: instruction <= 16'h0000;
		10'h20F: instruction <= 16'h0000;
		10'h210: instruction <= 16'h0000;
		10'h211: instruction <= 16'h0000;
		10'h212: instruction <= 16'h0000;
		10'h213: instruction <= 16'h0000;
		10'h214: instruction <= 16'h0000;
		10'h215: instruction <= 16'h0000;
		10'h216: instruction <= 16'h0000;
		10'h217: instruction <= 16'h0000;
		10'h218: instruction <= 16'h0000;
		10'h219: instruction <= 16'h0000;
		10'h21A: instruction <= 16'h0000;
		10'h21B: instruction <= 16'h0000;
		10'h21C: instruction <= 16'h0000;
		10'h21D: instruction <= 16'h0000;
		10'h21E: instruction <= 16'h0000;
		10'h21F: instruction <= 16'h0000;
		10'h220: instruction <= 16'h0000;
		10'h221: instruction <= 16'h0000;
		10'h222: instruction <= 16'h0000;
		10'h223: instruction <= 16'h0000;
		10'h224: instruction <= 16'h0000;
		10'h225: instruction <= 16'h0000;
		10'h226: instruction <= 16'h0000;
		10'h227: instruction <= 16'h0000;
		10'h228: instruction <= 16'h0000;
		10'h229: instruction <= 16'h0000;
		10'h22A: instruction <= 16'h0000;
		10'h22B: instruction <= 16'h0000;
		10'h22C: instruction <= 16'h0000;
		10'h22D: instruction <= 16'h0000;
		10'h22E: instruction <= 16'h0000;
		10'h22F: instruction <= 16'h0000;
		10'h230: instruction <= 16'h0000;
		10'h231: instruction <= 16'h0000;
		10'h232: instruction <= 16'h0000;
		10'h233: instruction <= 16'h0000;
		10'h234: instruction <= 16'h0000;
		10'h235: instruction <= 16'h0000;
		10'h236: instruction <= 16'h0000;
		10'h237: instruction <= 16'h0000;
		10'h238: instruction <= 16'h0000;
		10'h239: instruction <= 16'h0000;
		10'h23A: instruction <= 16'h0000;
		10'h23B: instruction <= 16'h0000;
		10'h23C: instruction <= 16'h0000;
		10'h23D: instruction <= 16'h0000;
		10'h23E: instruction <= 16'h0000;
		10'h23F: instruction <= 16'h0000;
		10'h240: instruction <= 16'h0000;
		10'h241: instruction <= 16'h0000;
		10'h242: instruction <= 16'h0000;
		10'h243: instruction <= 16'h0000;
		10'h244: instruction <= 16'h0000;
		10'h245: instruction <= 16'h0000;
		10'h246: instruction <= 16'h0000;
		10'h247: instruction <= 16'h0000;
		10'h248: instruction <= 16'h0000;
		10'h249: instruction <= 16'h0000;
		10'h24A: instruction <= 16'h0000;
		10'h24B: instruction <= 16'h0000;
		10'h24C: instruction <= 16'h0000;
		10'h24D: instruction <= 16'h0000;
		10'h24E: instruction <= 16'h0000;
		10'h24F: instruction <= 16'h0000;
		10'h250: instruction <= 16'h0000;
		10'h251: instruction <= 16'h0000;
		10'h252: instruction <= 16'h0000;
		10'h253: instruction <= 16'h0000;
		10'h254: instruction <= 16'h0000;
		10'h255: instruction <= 16'h0000;
		10'h256: instruction <= 16'h0000;
		10'h257: instruction <= 16'h0000;
		10'h258: instruction <= 16'h0000;
		10'h259: instruction <= 16'h0000;
		10'h25A: instruction <= 16'h0000;
		10'h25B: instruction <= 16'h0000;
		10'h25C: instruction <= 16'h0000;
		10'h25D: instruction <= 16'h0000;
		10'h25E: instruction <= 16'h0000;
		10'h25F: instruction <= 16'h0000;
		10'h260: instruction <= 16'h0000;
		10'h261: instruction <= 16'h0000;
		10'h262: instruction <= 16'h0000;
		10'h263: instruction <= 16'h0000;
		10'h264: instruction <= 16'h0000;
		10'h265: instruction <= 16'h0000;
		10'h266: instruction <= 16'h0000;
		10'h267: instruction <= 16'h0000;
		10'h268: instruction <= 16'h0000;
		10'h269: instruction <= 16'h0000;
		10'h26A: instruction <= 16'h0000;
		10'h26B: instruction <= 16'h0000;
		10'h26C: instruction <= 16'h0000;
		10'h26D: instruction <= 16'h0000;
		10'h26E: instruction <= 16'h0000;
		10'h26F: instruction <= 16'h0000;
		10'h270: instruction <= 16'h0000;
		10'h271: instruction <= 16'h0000;
		10'h272: instruction <= 16'h0000;
		10'h273: instruction <= 16'h0000;
		10'h274: instruction <= 16'h0000;
		10'h275: instruction <= 16'h0000;
		10'h276: instruction <= 16'h0000;
		10'h277: instruction <= 16'h0000;
		10'h278: instruction <= 16'h0000;
		10'h279: instruction <= 16'h0000;
		10'h27A: instruction <= 16'h0000;
		10'h27B: instruction <= 16'h0000;
		10'h27C: instruction <= 16'h0000;
		10'h27D: instruction <= 16'h0000;
		10'h27E: instruction <= 16'h0000;
		10'h27F: instruction <= 16'h0000;
		10'h280: instruction <= 16'h0000;
		10'h281: instruction <= 16'h0000;
		10'h282: instruction <= 16'h0000;
		10'h283: instruction <= 16'h0000;
		10'h284: instruction <= 16'h0000;
		10'h285: instruction <= 16'h0000;
		10'h286: instruction <= 16'h0000;
		10'h287: instruction <= 16'h0000;
		10'h288: instruction <= 16'h0000;
		10'h289: instruction <= 16'h0000;
		10'h28A: instruction <= 16'h0000;
		10'h28B: instruction <= 16'h0000;
		10'h28C: instruction <= 16'h0000;
		10'h28D: instruction <= 16'h0000;
		10'h28E: instruction <= 16'h0000;
		10'h28F: instruction <= 16'h0000;
		10'h290: instruction <= 16'h0000;
		10'h291: instruction <= 16'h0000;
		10'h292: instruction <= 16'h0000;
		10'h293: instruction <= 16'h0000;
		10'h294: instruction <= 16'h0000;
		10'h295: instruction <= 16'h0000;
		10'h296: instruction <= 16'h0000;
		10'h297: instruction <= 16'h0000;
		10'h298: instruction <= 16'h0000;
		10'h299: instruction <= 16'h0000;
		10'h29A: instruction <= 16'h0000;
		10'h29B: instruction <= 16'h0000;
		10'h29C: instruction <= 16'h0000;
		10'h29D: instruction <= 16'h0000;
		10'h29E: instruction <= 16'h0000;
		10'h29F: instruction <= 16'h0000;
		10'h2A0: instruction <= 16'h0000;
		10'h2A1: instruction <= 16'h0000;
		10'h2A2: instruction <= 16'h0000;
		10'h2A3: instruction <= 16'h0000;
		10'h2A4: instruction <= 16'h0000;
		10'h2A5: instruction <= 16'h0000;
		10'h2A6: instruction <= 16'h0000;
		10'h2A7: instruction <= 16'h0000;
		10'h2A8: instruction <= 16'h0000;
		10'h2A9: instruction <= 16'h0000;
		10'h2AA: instruction <= 16'h0000;
		10'h2AB: instruction <= 16'h0000;
		10'h2AC: instruction <= 16'h0000;
		10'h2AD: instruction <= 16'h0000;
		10'h2AE: instruction <= 16'h0000;
		10'h2AF: instruction <= 16'h0000;
		10'h2B0: instruction <= 16'h0000;
		10'h2B1: instruction <= 16'h0000;
		10'h2B2: instruction <= 16'h0000;
		10'h2B3: instruction <= 16'h0000;
		10'h2B4: instruction <= 16'h0000;
		10'h2B5: instruction <= 16'h0000;
		10'h2B6: instruction <= 16'h0000;
		10'h2B7: instruction <= 16'h0000;
		10'h2B8: instruction <= 16'h0000;
		10'h2B9: instruction <= 16'h0000;
		10'h2BA: instruction <= 16'h0000;
		10'h2BB: instruction <= 16'h0000;
		10'h2BC: instruction <= 16'h0000;
		10'h2BD: instruction <= 16'h0000;
		10'h2BE: instruction <= 16'h0000;
		10'h2BF: instruction <= 16'h0000;
		10'h2C0: instruction <= 16'h0000;
		10'h2C1: instruction <= 16'h0000;
		10'h2C2: instruction <= 16'h0000;
		10'h2C3: instruction <= 16'h0000;
		10'h2C4: instruction <= 16'h0000;
		10'h2C5: instruction <= 16'h0000;
		10'h2C6: instruction <= 16'h0000;
		10'h2C7: instruction <= 16'h0000;
		10'h2C8: instruction <= 16'h0000;
		10'h2C9: instruction <= 16'h0000;
		10'h2CA: instruction <= 16'h0000;
		10'h2CB: instruction <= 16'h0000;
		10'h2CC: instruction <= 16'h0000;
		10'h2CD: instruction <= 16'h0000;
		10'h2CE: instruction <= 16'h0000;
		10'h2CF: instruction <= 16'h0000;
		10'h2D0: instruction <= 16'h0000;
		10'h2D1: instruction <= 16'h0000;
		10'h2D2: instruction <= 16'h0000;
		10'h2D3: instruction <= 16'h0000;
		10'h2D4: instruction <= 16'h0000;
		10'h2D5: instruction <= 16'h0000;
		10'h2D6: instruction <= 16'h0000;
		10'h2D7: instruction <= 16'h0000;
		10'h2D8: instruction <= 16'h0000;
		10'h2D9: instruction <= 16'h0000;
		10'h2DA: instruction <= 16'h0000;
		10'h2DB: instruction <= 16'h0000;
		10'h2DC: instruction <= 16'h0000;
		10'h2DD: instruction <= 16'h0000;
		10'h2DE: instruction <= 16'h0000;
		10'h2DF: instruction <= 16'h0000;
		10'h2E0: instruction <= 16'h0000;
		10'h2E1: instruction <= 16'h0000;
		10'h2E2: instruction <= 16'h0000;
		10'h2E3: instruction <= 16'h0000;
		10'h2E4: instruction <= 16'h0000;
		10'h2E5: instruction <= 16'h0000;
		10'h2E6: instruction <= 16'h0000;
		10'h2E7: instruction <= 16'h0000;
		10'h2E8: instruction <= 16'h0000;
		10'h2E9: instruction <= 16'h0000;
		10'h2EA: instruction <= 16'h0000;
		10'h2EB: instruction <= 16'h0000;
		10'h2EC: instruction <= 16'h0000;
		10'h2ED: instruction <= 16'h0000;
		10'h2EE: instruction <= 16'h0000;
		10'h2EF: instruction <= 16'h0000;
		10'h2F0: instruction <= 16'h0000;
		10'h2F1: instruction <= 16'h0000;
		10'h2F2: instruction <= 16'h0000;
		10'h2F3: instruction <= 16'h0000;
		10'h2F4: instruction <= 16'h0000;
		10'h2F5: instruction <= 16'h0000;
		10'h2F6: instruction <= 16'h0000;
		10'h2F7: instruction <= 16'h0000;
		10'h2F8: instruction <= 16'h0000;
		10'h2F9: instruction <= 16'h0000;
		10'h2FA: instruction <= 16'h0000;
		10'h2FB: instruction <= 16'h0000;
		10'h2FC: instruction <= 16'h0000;
		10'h2FD: instruction <= 16'h0000;
		10'h2FE: instruction <= 16'h0000;
		10'h2FF: instruction <= 16'h0000;
		10'h300: instruction <= 16'h0000;
		10'h301: instruction <= 16'h0000;
		10'h302: instruction <= 16'h0000;
		10'h303: instruction <= 16'h0000;
		10'h304: instruction <= 16'h0000;
		10'h305: instruction <= 16'h0000;
		10'h306: instruction <= 16'h0000;
		10'h307: instruction <= 16'h0000;
		10'h308: instruction <= 16'h0000;
		10'h309: instruction <= 16'h0000;
		10'h30A: instruction <= 16'h0000;
		10'h30B: instruction <= 16'h0000;
		10'h30C: instruction <= 16'h0000;
		10'h30D: instruction <= 16'h0000;
		10'h30E: instruction <= 16'h0000;
		10'h30F: instruction <= 16'h0000;
		10'h310: instruction <= 16'h0000;
		10'h311: instruction <= 16'h0000;
		10'h312: instruction <= 16'h0000;
		10'h313: instruction <= 16'h0000;
		10'h314: instruction <= 16'h0000;
		10'h315: instruction <= 16'h0000;
		10'h316: instruction <= 16'h0000;
		10'h317: instruction <= 16'h0000;
		10'h318: instruction <= 16'h0000;
		10'h319: instruction <= 16'h0000;
		10'h31A: instruction <= 16'h0000;
		10'h31B: instruction <= 16'h0000;
		10'h31C: instruction <= 16'h0000;
		10'h31D: instruction <= 16'h0000;
		10'h31E: instruction <= 16'h0000;
		10'h31F: instruction <= 16'h0000;
		10'h320: instruction <= 16'h0000;
		10'h321: instruction <= 16'h0000;
		10'h322: instruction <= 16'h0000;
		10'h323: instruction <= 16'h0000;
		10'h324: instruction <= 16'h0000;
		10'h325: instruction <= 16'h0000;
		10'h326: instruction <= 16'h0000;
		10'h327: instruction <= 16'h0000;
		10'h328: instruction <= 16'h0000;
		10'h329: instruction <= 16'h0000;
		10'h32A: instruction <= 16'h0000;
		10'h32B: instruction <= 16'h0000;
		10'h32C: instruction <= 16'h0000;
		10'h32D: instruction <= 16'h0000;
		10'h32E: instruction <= 16'h0000;
		10'h32F: instruction <= 16'h0000;
		10'h330: instruction <= 16'h0000;
		10'h331: instruction <= 16'h0000;
		10'h332: instruction <= 16'h0000;
		10'h333: instruction <= 16'h0000;
		10'h334: instruction <= 16'h0000;
		10'h335: instruction <= 16'h0000;
		10'h336: instruction <= 16'h0000;
		10'h337: instruction <= 16'h0000;
		10'h338: instruction <= 16'h0000;
		10'h339: instruction <= 16'h0000;
		10'h33A: instruction <= 16'h0000;
		10'h33B: instruction <= 16'h0000;
		10'h33C: instruction <= 16'h0000;
		10'h33D: instruction <= 16'h0000;
		10'h33E: instruction <= 16'h0000;
		10'h33F: instruction <= 16'h0000;
		10'h340: instruction <= 16'h0000;
		10'h341: instruction <= 16'h0000;
		10'h342: instruction <= 16'h0000;
		10'h343: instruction <= 16'h0000;
		10'h344: instruction <= 16'h0000;
		10'h345: instruction <= 16'h0000;
		10'h346: instruction <= 16'h0000;
		10'h347: instruction <= 16'h0000;
		10'h348: instruction <= 16'h0000;
		10'h349: instruction <= 16'h0000;
		10'h34A: instruction <= 16'h0000;
		10'h34B: instruction <= 16'h0000;
		10'h34C: instruction <= 16'h0000;
		10'h34D: instruction <= 16'h0000;
		10'h34E: instruction <= 16'h0000;
		10'h34F: instruction <= 16'h0000;
		10'h350: instruction <= 16'h0000;
		10'h351: instruction <= 16'h0000;
		10'h352: instruction <= 16'h0000;
		10'h353: instruction <= 16'h0000;
		10'h354: instruction <= 16'h0000;
		10'h355: instruction <= 16'h0000;
		10'h356: instruction <= 16'h0000;
		10'h357: instruction <= 16'h0000;
		10'h358: instruction <= 16'h0000;
		10'h359: instruction <= 16'h0000;
		10'h35A: instruction <= 16'h0000;
		10'h35B: instruction <= 16'h0000;
		10'h35C: instruction <= 16'h0000;
		10'h35D: instruction <= 16'h0000;
		10'h35E: instruction <= 16'h0000;
		10'h35F: instruction <= 16'h0000;
		10'h360: instruction <= 16'h0000;
		10'h361: instruction <= 16'h0000;
		10'h362: instruction <= 16'h0000;
		10'h363: instruction <= 16'h0000;
		10'h364: instruction <= 16'h0000;
		10'h365: instruction <= 16'h0000;
		10'h366: instruction <= 16'h0000;
		10'h367: instruction <= 16'h0000;
		10'h368: instruction <= 16'h0000;
		10'h369: instruction <= 16'h0000;
		10'h36A: instruction <= 16'h0000;
		10'h36B: instruction <= 16'h0000;
		10'h36C: instruction <= 16'h0000;
		10'h36D: instruction <= 16'h0000;
		10'h36E: instruction <= 16'h0000;
		10'h36F: instruction <= 16'h0000;
		10'h370: instruction <= 16'h0000;
		10'h371: instruction <= 16'h0000;
		10'h372: instruction <= 16'h0000;
		10'h373: instruction <= 16'h0000;
		10'h374: instruction <= 16'h0000;
		10'h375: instruction <= 16'h0000;
		10'h376: instruction <= 16'h0000;
		10'h377: instruction <= 16'h0000;
		10'h378: instruction <= 16'h0000;
		10'h379: instruction <= 16'h0000;
		10'h37A: instruction <= 16'h0000;
		10'h37B: instruction <= 16'h0000;
		10'h37C: instruction <= 16'h0000;
		10'h37D: instruction <= 16'h0000;
		10'h37E: instruction <= 16'h0000;
		10'h37F: instruction <= 16'h0000;
		10'h380: instruction <= 16'h0000;
		10'h381: instruction <= 16'h0000;
		10'h382: instruction <= 16'h0000;
		10'h383: instruction <= 16'h0000;
		10'h384: instruction <= 16'h0000;
		10'h385: instruction <= 16'h0000;
		10'h386: instruction <= 16'h0000;
		10'h387: instruction <= 16'h0000;
		10'h388: instruction <= 16'h0000;
		10'h389: instruction <= 16'h0000;
		10'h38A: instruction <= 16'h0000;
		10'h38B: instruction <= 16'h0000;
		10'h38C: instruction <= 16'h0000;
		10'h38D: instruction <= 16'h0000;
		10'h38E: instruction <= 16'h0000;
		10'h38F: instruction <= 16'h0000;
		10'h390: instruction <= 16'h0000;
		10'h391: instruction <= 16'h0000;
		10'h392: instruction <= 16'h0000;
		10'h393: instruction <= 16'h0000;
		10'h394: instruction <= 16'h0000;
		10'h395: instruction <= 16'h0000;
		10'h396: instruction <= 16'h0000;
		10'h397: instruction <= 16'h0000;
		10'h398: instruction <= 16'h0000;
		10'h399: instruction <= 16'h0000;
		10'h39A: instruction <= 16'h0000;
		10'h39B: instruction <= 16'h0000;
		10'h39C: instruction <= 16'h0000;
		10'h39D: instruction <= 16'h0000;
		10'h39E: instruction <= 16'h0000;
		10'h39F: instruction <= 16'h0000;
		10'h3A0: instruction <= 16'h0000;
		10'h3A1: instruction <= 16'h0000;
		10'h3A2: instruction <= 16'h0000;
		10'h3A3: instruction <= 16'h0000;
		10'h3A4: instruction <= 16'h0000;
		10'h3A5: instruction <= 16'h0000;
		10'h3A6: instruction <= 16'h0000;
		10'h3A7: instruction <= 16'h0000;
		10'h3A8: instruction <= 16'h0000;
		10'h3A9: instruction <= 16'h0000;
		10'h3AA: instruction <= 16'h0000;
		10'h3AB: instruction <= 16'h0000;
		10'h3AC: instruction <= 16'h0000;
		10'h3AD: instruction <= 16'h0000;
		10'h3AE: instruction <= 16'h0000;
		10'h3AF: instruction <= 16'h0000;
		10'h3B0: instruction <= 16'h0000;
		10'h3B1: instruction <= 16'h0000;
		10'h3B2: instruction <= 16'h0000;
		10'h3B3: instruction <= 16'h0000;
		10'h3B4: instruction <= 16'h0000;
		10'h3B5: instruction <= 16'h0000;
		10'h3B6: instruction <= 16'h0000;
		10'h3B7: instruction <= 16'h0000;
		10'h3B8: instruction <= 16'h0000;
		10'h3B9: instruction <= 16'h0000;
		10'h3BA: instruction <= 16'h0000;
		10'h3BB: instruction <= 16'h0000;
		10'h3BC: instruction <= 16'h0000;
		10'h3BD: instruction <= 16'h0000;
		10'h3BE: instruction <= 16'h0000;
		10'h3BF: instruction <= 16'h0000;
		10'h3C0: instruction <= 16'h0000;
		10'h3C1: instruction <= 16'h0000;
		10'h3C2: instruction <= 16'h0000;
		10'h3C3: instruction <= 16'h0000;
		10'h3C4: instruction <= 16'h0000;
		10'h3C5: instruction <= 16'h0000;
		10'h3C6: instruction <= 16'h0000;
		10'h3C7: instruction <= 16'h0000;
		10'h3C8: instruction <= 16'h0000;
		10'h3C9: instruction <= 16'h0000;
		10'h3CA: instruction <= 16'h0000;
		10'h3CB: instruction <= 16'h0000;
		10'h3CC: instruction <= 16'h0000;
		10'h3CD: instruction <= 16'h0000;
		10'h3CE: instruction <= 16'h0000;
		10'h3CF: instruction <= 16'h0000;
		10'h3D0: instruction <= 16'h0000;
		10'h3D1: instruction <= 16'h0000;
		10'h3D2: instruction <= 16'h0000;
		10'h3D3: instruction <= 16'h0000;
		10'h3D4: instruction <= 16'h0000;
		10'h3D5: instruction <= 16'h0000;
		10'h3D6: instruction <= 16'h0000;
		10'h3D7: instruction <= 16'h0000;
		10'h3D8: instruction <= 16'h0000;
		10'h3D9: instruction <= 16'h0000;
		10'h3DA: instruction <= 16'h0000;
		10'h3DB: instruction <= 16'h0000;
		10'h3DC: instruction <= 16'h0000;
		10'h3DD: instruction <= 16'h0000;
		10'h3DE: instruction <= 16'h0000;
		10'h3DF: instruction <= 16'h0000;
		10'h3E0: instruction <= 16'h0000;
		10'h3E1: instruction <= 16'h0000;
		10'h3E2: instruction <= 16'h0000;
		10'h3E3: instruction <= 16'h0000;
		10'h3E4: instruction <= 16'h0000;
		10'h3E5: instruction <= 16'h0000;
		10'h3E6: instruction <= 16'h0000;
		10'h3E7: instruction <= 16'h0000;
		10'h3E8: instruction <= 16'h0000;
		10'h3E9: instruction <= 16'h0000;
		10'h3EA: instruction <= 16'h0000;
		10'h3EB: instruction <= 16'h0000;
		10'h3EC: instruction <= 16'h0000;
		10'h3ED: instruction <= 16'h0000;
		10'h3EE: instruction <= 16'h0000;
		10'h3EF: instruction <= 16'h0000;
		10'h3F0: instruction <= 16'h0000;
		10'h3F1: instruction <= 16'h0000;
		10'h3F2: instruction <= 16'h0000;
		10'h3F3: instruction <= 16'h0000;
		10'h3F4: instruction <= 16'h0000;
		10'h3F5: instruction <= 16'h0000;
		10'h3F6: instruction <= 16'h0000;
		10'h3F7: instruction <= 16'h0000;
		10'h3F8: instruction <= 16'h0000;
		10'h3F9: instruction <= 16'h0000;
		10'h3FA: instruction <= 16'h0000;
		10'h3FB: instruction <= 16'h0000;
		10'h3FC: instruction <= 16'h0000;
		10'h3FD: instruction <= 16'h0000;
		10'h3FE: instruction <= 16'h0000;
		10'h3FF: instruction <= 16'h0000;
		default: instruction <= 16'h0000;
	endcase
end
endmodule
